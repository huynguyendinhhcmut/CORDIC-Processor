module multiply32x32 (
	input wire [31:0] a, b,
	output wire [63:0] mul
);

wire [31:0] sum1,  sum2,  sum3,  sum4,  sum5,  sum6,  sum7,  sum8,  sum9,  sum10,
       	    sum11, sum12, sum13, sum14, sum15, sum16, sum17, sum18, sum19, sum20, 
	    sum21, sum22, sum23, sum24, sum25, sum26, sum27, sum28, sum29, sum30, sum31;
wire carry1,  carry2,  carry3,  carry4,  carry5,  carry6,  carry7,  carry8,  carry9,  carry10, 
     carry11, carry12, carry13, carry14, carry15, carry16, carry17, carry18, carry19, carry20, 
     carry21, carry22, carry23, carry24, carry25, carry26, carry27, carry28, carry29, carry30, carry31;

and (mul[0], a[0], b[0]);

fullAdder32b fa1 (.sum(sum1), .a0(a[1] & b[0]),   .a1(a[2] & b[0]),   .a2(a[3] & b[0]),   .a3(a[4] & b[0]),   .a4(a[5] & b[0]),   .a5(a[6] & b[0]),   .a6(a[7] & b[0]),   .a7(a[8] & b[0]),
			      .a8(a[9] & b[0]),   .a9(a[10] & b[0]),  .a10(a[11] & b[0]), .a11(a[12] & b[0]), .a12(a[13] & b[0]), .a13(a[14] & b[0]), .a14(a[15] & b[0]), .a15(a[16] & b[0]),
			      .a16(a[9] & b[0]),  .a17(a[10] & b[0]), .a18(a[11] & b[0]), .a19(a[12] & b[0]), .a20(a[13] & b[0]), .a21(a[14] & b[0]), .a22(a[15] & b[0]), .a23(a[16] & b[0]),
	                      .a24(a[25] & b[0]), .a25(a[26] & b[0]), .a26(a[27] & b[0]), .a27(a[28] & b[0]), .a28(a[29] & b[0]), .a29(a[30] & b[0]), .a30(a[31] & b[0]), .a31(1'b0),
			  
			      .b0(a[0] & b[1]),   .b1(a[1] & b[1]),   .b2(a[2] & b[1]),   .b3(a[3] & b[1]),   .b4(a[4] & b[1]),   .b5(a[5] & b[1]),   .b6(a[6] & b[1]),   .b7(a[7] & b[1]),
			      .b8(a[8] & b[1]),   .b9(a[9] & b[1]),   .b10(a[10] & b[1]), .b11(a[12] & b[1]), .b12(a[12] & b[1]), .b13(a[13] & b[1]), .b14(a[14] & b[1]), .b15(a[15] & b[1]),
			      .b16(a[16] & b[1]), .b17(a[17] & b[1]), .b18(a[18] & b[1]), .b19(a[19] & b[1]), .b20(a[20] & b[1]), .b21(a[21] & b[1]), .b22(a[22] & b[1]), .b23(a[23] & b[1]),
	                      .b24(a[24] & b[1]), .b25(a[25] & b[1]), .b26(a[26] & b[1]), .b27(a[27] & b[1]), .b28(a[28] & b[1]), .b29(a[29] & b[1]), .b30(a[30] & b[1]), .b31(a[31] & b[1]),	  
	          .cin(1'b0), .cout(carry1));

fullAdder32b fa2 (.sum(sum2), .a0(sum1[1]),   .a1(sum1[2]),   .a2(sum1[3]),   .a3(sum1[4]),   .a4(sum1[5]),   .a5(sum1[6]),   .a6(sum1[7]),   .a7(sum1[8]),   .a8(sum1[9]),   .a9(sum1[10]),  .a10(sum1[11]), 
		              .a11(sum1[12]), .a12(sum1[13]), .a13(sum1[14]), .a14(sum1[15]), .a15(sum1[16]), .a16(sum1[17]), .a17(sum1[18]), .a18(sum1[19]), .a19(sum1[20]), .a20(sum1[21]), .a21(sum1[22]),
			      .a22(sum1[23]), .a23(sum1[24]), .a24(sum1[25]), .a25(sum1[26]), .a26(sum1[27]), .a27(sum1[28]), .a28(sum1[29]), .a29(sum1[30]), .a30(sum1[31]), .a31(carry1), 

			      .b0(a[0] & b[2]),   .b1(a[1] & b[2]),   .b2(a[2] & b[2]),   .b3(a[3] & b[2]),   .b4(a[4] & b[2]),   .b5(a[5] & b[2]),   .b6(a[6] & b[2]),   .b7(a[7] & b[2]),
			      .b8(a[8] & b[2]),   .b9(a[9] & b[2]),   .b10(a[10] & b[2]), .b11(a[12] & b[2]), .b12(a[12] & b[2]), .b13(a[13] & b[2]), .b14(a[14] & b[2]), .b15(a[15] & b[2]),
			      .b16(a[16] & b[2]), .b17(a[17] & b[2]), .b18(a[18] & b[2]), .b19(a[19] & b[2]), .b20(a[20] & b[2]), .b21(a[21] & b[2]), .b22(a[22] & b[2]), .b23(a[23] & b[2]),
	                      .b24(a[24] & b[2]), .b25(a[25] & b[2]), .b26(a[26] & b[2]), .b27(a[27] & b[2]), .b28(a[28] & b[2]), .b29(a[29] & b[2]), .b30(a[30] & b[2]), .b31(a[31] & b[2]),	  
	          .cin(1'b0), .cout(carry2));


fullAdder32b fa3 (.sum(sum3), .a0(sum2[1]),   .a1(sum2[2]),   .a2(sum2[3]),   .a3(sum2[4]),   .a4(sum2[5]),   .a5(sum2[6]),   .a6(sum2[7]),   .a7(sum2[8]),   .a8(sum2[9]),   .a9(sum2[10]),  .a10(sum2[11]), 
		              .a11(sum2[12]), .a12(sum2[13]), .a13(sum2[14]), .a14(sum2[15]), .a15(sum2[16]), .a16(sum2[17]), .a17(sum2[18]), .a18(sum2[19]), .a19(sum2[20]), .a20(sum2[21]), .a21(sum2[22]),
			      .a22(sum2[23]), .a23(sum2[24]), .a24(sum2[25]), .a25(sum2[26]), .a26(sum2[27]), .a27(sum2[28]), .a28(sum2[29]), .a29(sum2[30]), .a30(sum2[31]), .a31(carry2), 

			      .b0(a[0] & b[3]),   .b1(a[1] & b[3]),   .b2(a[2] & b[3]),   .b3(a[3] & b[3]),   .b4(a[4] & b[3]),   .b5(a[5] & b[3]),   .b6(a[6] & b[3]),   .b7(a[7] & b[3]),
			      .b8(a[8] & b[3]),   .b9(a[9] & b[3]),   .b10(a[10] & b[3]), .b11(a[12] & b[3]), .b12(a[12] & b[3]), .b13(a[13] & b[3]), .b14(a[14] & b[3]), .b15(a[15] & b[3]),
			      .b16(a[16] & b[3]), .b17(a[17] & b[3]), .b18(a[18] & b[3]), .b19(a[19] & b[3]), .b20(a[20] & b[3]), .b21(a[21] & b[3]), .b22(a[22] & b[3]), .b23(a[23] & b[3]),
	                      .b24(a[24] & b[3]), .b25(a[25] & b[3]), .b26(a[26] & b[3]), .b27(a[27] & b[3]), .b28(a[28] & b[3]), .b29(a[29] & b[3]), .b30(a[30] & b[3]), .b31(a[31] & b[3]),	  
	          .cin(1'b0), .cout(carry3));

fullAdder32b fa4 (.sum(sum4), .a0(sum3[1]),   .a1(sum3[2]),   .a2(sum3[3]),   .a3(sum3[4]),   .a4(sum3[5]),   .a5(sum3[6]),   .a6(sum3[7]),   .a7(sum3[8]),   .a8(sum3[9]),   .a9(sum3[10]),  .a10(sum3[11]), 
		              .a11(sum3[12]), .a12(sum3[13]), .a13(sum3[14]), .a14(sum3[15]), .a15(sum3[16]), .a16(sum3[17]), .a17(sum3[18]), .a18(sum3[19]), .a19(sum3[20]), .a20(sum3[21]), .a21(sum3[22]),
			      .a22(sum3[23]), .a23(sum3[24]), .a24(sum3[25]), .a25(sum3[26]), .a26(sum3[27]), .a27(sum3[28]), .a28(sum3[29]), .a29(sum3[30]), .a30(sum3[31]), .a31(carry3), 

			      .b0(a[0] & b[4]),   .b1(a[1] & b[4]),   .b2(a[2] & b[4]),   .b3(a[3] & b[4]),   .b4(a[4] & b[4]),   .b5(a[5] & b[4]),   .b6(a[6] & b[4]),   .b7(a[7] & b[4]),
			      .b8(a[8] & b[4]),   .b9(a[9] & b[4]),   .b10(a[10] & b[4]), .b11(a[12] & b[4]), .b12(a[12] & b[4]), .b13(a[13] & b[4]), .b14(a[14] & b[4]), .b15(a[15] & b[4]),
			      .b16(a[16] & b[4]), .b17(a[17] & b[4]), .b18(a[18] & b[4]), .b19(a[19] & b[4]), .b20(a[20] & b[4]), .b21(a[21] & b[4]), .b22(a[22] & b[4]), .b23(a[23] & b[4]),
	                      .b24(a[24] & b[4]), .b25(a[25] & b[4]), .b26(a[26] & b[4]), .b27(a[27] & b[4]), .b28(a[28] & b[4]), .b29(a[29] & b[4]), .b30(a[30] & b[4]), .b31(a[31] & b[4]),	  
	          .cin(1'b0), .cout(carry4));

fullAdder32b fa5 (.sum(sum5), .a0(sum4[1]),   .a1(sum4[2]),   .a2(sum4[3]),   .a3(sum4[4]),   .a4(sum4[5]),   .a5(sum4[6]),   .a6(sum4[7]),   .a7(sum4[8]),   .a8(sum4[9]),   .a9(sum4[10]),  .a10(sum4[11]), 
		              .a11(sum4[12]), .a12(sum4[13]), .a13(sum4[14]), .a14(sum4[15]), .a15(sum4[16]), .a16(sum4[17]), .a17(sum4[18]), .a18(sum4[19]), .a19(sum4[20]), .a20(sum4[21]), .a21(sum4[22]),
			      .a22(sum4[23]), .a23(sum4[24]), .a24(sum4[25]), .a25(sum4[26]), .a26(sum4[27]), .a27(sum4[28]), .a28(sum4[29]), .a29(sum4[30]), .a30(sum4[31]), .a31(carry4), 

			      .b0(a[0] & b[5]),   .b1(a[1] & b[5]),   .b2(a[2] & b[5]),   .b3(a[3] & b[5]),   .b4(a[4] & b[5]),   .b5(a[5] & b[5]),   .b6(a[6] & b[5]),   .b7(a[7] & b[5]),
			      .b8(a[8] & b[5]),   .b9(a[9] & b[5]),   .b10(a[10] & b[5]), .b11(a[12] & b[5]), .b12(a[12] & b[5]), .b13(a[13] & b[5]), .b14(a[14] & b[5]), .b15(a[15] & b[5]),
			      .b16(a[16] & b[5]), .b17(a[17] & b[5]), .b18(a[18] & b[5]), .b19(a[19] & b[5]), .b20(a[20] & b[5]), .b21(a[21] & b[5]), .b22(a[22] & b[5]), .b23(a[23] & b[5]),
	                      .b24(a[24] & b[5]), .b25(a[25] & b[5]), .b26(a[26] & b[5]), .b27(a[27] & b[5]), .b28(a[28] & b[5]), .b29(a[29] & b[5]), .b30(a[30] & b[5]), .b31(a[31] & b[5]),	  
	          .cin(1'b0), .cout(carry5));

fullAdder32b fa6 (.sum(sum6), .a0(sum5[1]),   .a1(sum5[2]),   .a2(sum5[3]),   .a3(sum5[4]),   .a4(sum5[5]),   .a5(sum5[6]),   .a6(sum5[7]),   .a7(sum5[8]),   .a8(sum5[9]),   .a9(sum5[10]),  .a10(sum5[11]), 
		              .a11(sum5[12]), .a12(sum5[13]), .a13(sum5[14]), .a14(sum5[15]), .a15(sum5[16]), .a16(sum5[17]), .a17(sum5[18]), .a18(sum5[19]), .a19(sum5[20]), .a20(sum5[21]), .a21(sum5[22]),
			      .a22(sum5[23]), .a23(sum5[24]), .a24(sum5[25]), .a25(sum5[26]), .a26(sum5[27]), .a27(sum5[28]), .a28(sum5[29]), .a29(sum5[30]), .a30(sum5[31]), .a31(carry5), 

			      .b0(a[0] & b[6]),   .b1(a[1] & b[6]),   .b2(a[2] & b[6]),   .b3(a[3] & b[6]),   .b4(a[4] & b[6]),   .b5(a[5] & b[6]),   .b6(a[6] & b[6]),   .b7(a[7] & b[6]),
			      .b8(a[8] & b[6]),   .b9(a[9] & b[6]),   .b10(a[10] & b[6]), .b11(a[12] & b[6]), .b12(a[12] & b[6]), .b13(a[13] & b[6]), .b14(a[14] & b[6]), .b15(a[15] & b[6]),
			      .b16(a[16] & b[6]), .b17(a[17] & b[6]), .b18(a[18] & b[6]), .b19(a[19] & b[6]), .b20(a[20] & b[6]), .b21(a[21] & b[6]), .b22(a[22] & b[6]), .b23(a[23] & b[6]),
	                      .b24(a[24] & b[6]), .b25(a[25] & b[6]), .b26(a[26] & b[6]), .b27(a[27] & b[6]), .b28(a[28] & b[6]), .b29(a[29] & b[6]), .b30(a[30] & b[6]), .b31(a[31] & b[6]),	  
	          .cin(1'b0), .cout(carry6));

fullAdder32b fa7 (.sum(sum7), .a0(sum6[1]),   .a1(sum6[2]),   .a2(sum6[3]),   .a3(sum6[4]),   .a4(sum6[5]),   .a5(sum6[6]),   .a6(sum6[7]),   .a7(sum6[8]),   .a8(sum6[9]),   .a9(sum6[10]),  .a10(sum6[11]), 
		              .a11(sum6[12]), .a12(sum6[13]), .a13(sum6[14]), .a14(sum6[15]), .a15(sum6[16]), .a16(sum6[17]), .a17(sum6[18]), .a18(sum6[19]), .a19(sum6[20]), .a20(sum6[21]), .a21(sum6[22]),
			      .a22(sum6[23]), .a23(sum6[24]), .a24(sum6[25]), .a25(sum6[26]), .a26(sum6[27]), .a27(sum6[28]), .a28(sum6[29]), .a29(sum6[30]), .a30(sum6[31]), .a31(carry6), 

			      .b0(a[0] & b[7]),   .b1(a[1] & b[7]),   .b2(a[2] & b[7]),   .b3(a[3] & b[7]),   .b4(a[4] & b[7]),   .b5(a[5] & b[7]),   .b6(a[6] & b[7]),   .b7(a[7] & b[7]),
			      .b8(a[8] & b[7]),   .b9(a[9] & b[7]),   .b10(a[10] & b[7]), .b11(a[12] & b[7]), .b12(a[12] & b[7]), .b13(a[13] & b[7]), .b14(a[14] & b[7]), .b15(a[15] & b[7]),
			      .b16(a[16] & b[7]), .b17(a[17] & b[7]), .b18(a[18] & b[7]), .b19(a[19] & b[7]), .b20(a[20] & b[7]), .b21(a[21] & b[7]), .b22(a[22] & b[7]), .b23(a[23] & b[7]),
	                      .b24(a[24] & b[7]), .b25(a[25] & b[7]), .b26(a[26] & b[7]), .b27(a[27] & b[7]), .b28(a[28] & b[7]), .b29(a[29] & b[7]), .b30(a[30] & b[7]), .b31(a[31] & b[7]),	  
	          .cin(1'b0), .cout(carry7));

fullAdder32b fa8 (.sum(sum8), .a0(sum7[1]),   .a1(sum7[2]),   .a2(sum7[3]),   .a3(sum7[4]),   .a4(sum7[5]),   .a5(sum7[6]),   .a6(sum7[7]),   .a7(sum7[8]),   .a8(sum7[9]),   .a9(sum7[10]),  .a10(sum7[11]), 
		              .a11(sum7[12]), .a12(sum7[13]), .a13(sum7[14]), .a14(sum7[15]), .a15(sum7[16]), .a16(sum7[17]), .a17(sum7[18]), .a18(sum7[19]), .a19(sum7[20]), .a20(sum7[21]), .a21(sum7[22]),
			      .a22(sum7[23]), .a23(sum7[24]), .a24(sum7[25]), .a25(sum7[26]), .a26(sum7[27]), .a27(sum7[28]), .a28(sum7[29]), .a29(sum7[30]), .a30(sum7[31]), .a31(carry7), 

			      .b0(a[0] & b[8]),   .b1(a[1] & b[8]),   .b2(a[2] & b[8]),   .b3(a[3] & b[8]),   .b4(a[4] & b[8]),   .b5(a[5] & b[8]),   .b6(a[6] & b[8]),   .b7(a[7] & b[8]),
			      .b8(a[8] & b[8]),   .b9(a[9] & b[8]),   .b10(a[10] & b[8]), .b11(a[12] & b[8]), .b12(a[12] & b[8]), .b13(a[13] & b[8]), .b14(a[14] & b[8]), .b15(a[15] & b[8]),
			      .b16(a[16] & b[8]), .b17(a[17] & b[8]), .b18(a[18] & b[8]), .b19(a[19] & b[8]), .b20(a[20] & b[8]), .b21(a[21] & b[8]), .b22(a[22] & b[8]), .b23(a[23] & b[8]),
	                      .b24(a[24] & b[8]), .b25(a[25] & b[8]), .b26(a[26] & b[8]), .b27(a[27] & b[8]), .b28(a[28] & b[8]), .b29(a[29] & b[8]), .b30(a[30] & b[8]), .b31(a[31] & b[8]),	  
	          .cin(1'b0), .cout(carry8));

fullAdder32b fa9 (.sum(sum9), .a0(sum8[1]),   .a1(sum8[2]),   .a2(sum8[3]),   .a3(sum8[4]),   .a4(sum8[5]),   .a5(sum8[6]),   .a6(sum8[7]),   .a7(sum8[8]),   .a8(sum8[9]),   .a9(sum8[10]),  .a10(sum8[11]), 
		              .a11(sum8[12]), .a12(sum8[13]), .a13(sum8[14]), .a14(sum8[15]), .a15(sum8[16]), .a16(sum8[17]), .a17(sum8[18]), .a18(sum8[19]), .a19(sum8[20]), .a20(sum8[21]), .a21(sum8[22]),
			      .a22(sum8[23]), .a23(sum8[24]), .a24(sum8[25]), .a25(sum8[26]), .a26(sum8[27]), .a27(sum8[28]), .a28(sum8[29]), .a29(sum8[30]), .a30(sum8[31]), .a31(carry8), 

			      .b0(a[0] & b[9]),   .b1(a[1] & b[9]),   .b2(a[2] & b[9]),   .b3(a[3] & b[9]),   .b4(a[4] & b[9]),   .b5(a[5] & b[9]),   .b6(a[6] & b[9]),   .b7(a[7] & b[9]),
			      .b8(a[8] & b[9]),   .b9(a[9] & b[9]),   .b10(a[10] & b[9]), .b11(a[12] & b[9]), .b12(a[12] & b[9]), .b13(a[13] & b[9]), .b14(a[14] & b[9]), .b15(a[15] & b[9]),
			      .b16(a[16] & b[9]), .b17(a[17] & b[9]), .b18(a[18] & b[9]), .b19(a[19] & b[9]), .b20(a[20] & b[9]), .b21(a[21] & b[9]), .b22(a[22] & b[9]), .b23(a[23] & b[9]),
	                      .b24(a[24] & b[9]), .b25(a[25] & b[9]), .b26(a[26] & b[9]), .b27(a[27] & b[9]), .b28(a[28] & b[9]), .b29(a[29] & b[9]), .b30(a[30] & b[9]), .b31(a[31] & b[9]),	  
	          .cin(1'b0), .cout(carry9));

fullAdder32b fa10 (.sum(sum10), .a0(sum9[1]),   .a1(sum9[2]),   .a2(sum9[3]),   .a3(sum9[4]),   .a4(sum9[5]),   .a5(sum9[6]),   .a6(sum9[7]),   .a7(sum9[8]),   .a8(sum9[9]),   .a9(sum9[10]),  .a10(sum9[11]), 
		                .a11(sum9[12]), .a12(sum9[13]), .a13(sum9[14]), .a14(sum9[15]), .a15(sum9[16]), .a16(sum9[17]), .a17(sum9[18]), .a18(sum9[19]), .a19(sum9[20]), .a20(sum9[21]), .a21(sum9[22]),
			        .a22(sum9[23]), .a23(sum9[24]), .a24(sum9[25]), .a25(sum9[26]), .a26(sum9[27]), .a27(sum9[28]), .a28(sum9[29]), .a29(sum9[30]), .a30(sum9[31]), .a31(carry9), 

			        .b0(a[0] & b[10]),   .b1(a[1] & b[10]),   .b2(a[2] & b[10]),   .b3(a[3] & b[10]),   .b4(a[4] & b[10]),   .b5(a[5] & b[10]),   .b6(a[6] & b[10]),   .b7(a[7] & b[10]),
			        .b8(a[8] & b[10]),   .b9(a[9] & b[10]),   .b10(a[10] & b[10]), .b11(a[12] & b[10]), .b12(a[12] & b[10]), .b13(a[13] & b[10]), .b14(a[14] & b[10]), .b15(a[15] & b[10]),
			        .b16(a[16] & b[10]), .b17(a[17] & b[10]), .b18(a[18] & b[10]), .b19(a[19] & b[10]), .b20(a[20] & b[10]), .b21(a[21] & b[10]), .b22(a[22] & b[10]), .b23(a[23] & b[10]),
	                        .b24(a[24] & b[10]), .b25(a[25] & b[10]), .b26(a[26] & b[10]), .b27(a[27] & b[10]), .b28(a[28] & b[10]), .b29(a[29] & b[10]), .b30(a[30] & b[10]), .b31(a[31] & b[10]),	  
	          .cin(1'b0), .cout(carry10));

fullAdder32b fa11 (.sum(sum11), .a0(sum10[1]),   .a1(sum10[2]),   .a2(sum10[3]),   .a3(sum10[4]),   .a4(sum10[5]),   .a5(sum10[6]),   .a6(sum10[7]),   .a7(sum10[8]),   .a8(sum10[9]),   .a9(sum10[10]),  .a10(sum10[11]), 
		                .a11(sum10[12]), .a12(sum10[13]), .a13(sum10[14]), .a14(sum10[15]), .a15(sum10[16]), .a16(sum10[17]), .a17(sum10[18]), .a18(sum10[19]), .a19(sum10[20]), .a20(sum10[21]), .a21(sum10[22]),
			        .a22(sum10[23]), .a23(sum10[24]), .a24(sum10[25]), .a25(sum10[26]), .a26(sum10[27]), .a27(sum10[28]), .a28(sum10[29]), .a29(sum10[30]), .a30(sum10[31]), .a31(carry10), 

			        .b0(a[0] & b[11]),   .b1(a[1] & b[11]),   .b2(a[2] & b[11]),   .b3(a[3] & b[11]),   .b4(a[4] & b[11]),   .b5(a[5] & b[11]),   .b6(a[6] & b[11]),   .b7(a[7] & b[11]),
			        .b8(a[8] & b[11]),   .b9(a[9] & b[11]),   .b10(a[10] & b[11]), .b11(a[12] & b[11]), .b12(a[12] & b[11]), .b13(a[13] & b[11]), .b14(a[14] & b[11]), .b15(a[15] & b[11]),
			        .b16(a[16] & b[11]), .b17(a[17] & b[11]), .b18(a[18] & b[11]), .b19(a[19] & b[11]), .b20(a[20] & b[11]), .b21(a[21] & b[11]), .b22(a[22] & b[11]), .b23(a[23] & b[11]),
	                        .b24(a[24] & b[11]), .b25(a[25] & b[11]), .b26(a[26] & b[11]), .b27(a[27] & b[11]), .b28(a[28] & b[11]), .b29(a[29] & b[11]), .b30(a[30] & b[11]), .b31(a[31] & b[11]),	  
	          .cin(1'b0), .cout(carry11));

fullAdder32b fa12 (.sum(sum12), .a0(sum11[1]),   .a1(sum11[2]),   .a2(sum11[3]),   .a3(sum11[4]),   .a4(sum11[5]),   .a5(sum11[6]),   .a6(sum11[7]),   .a7(sum11[8]),   .a8(sum11[9]),   .a9(sum11[10]),  .a10(sum11[11]), 
		                .a11(sum11[12]), .a12(sum11[13]), .a13(sum11[14]), .a14(sum11[15]), .a15(sum11[16]), .a16(sum11[17]), .a17(sum11[18]), .a18(sum11[19]), .a19(sum11[20]), .a20(sum11[21]), .a21(sum11[22]),
			        .a22(sum11[23]), .a23(sum11[24]), .a24(sum11[25]), .a25(sum11[26]), .a26(sum11[27]), .a27(sum11[28]), .a28(sum11[29]), .a29(sum11[30]), .a30(sum11[31]), .a31(carry11), 

			        .b0(a[0] & b[12]),   .b1(a[1] & b[12]),   .b2(a[2] & b[12]),   .b3(a[3] & b[12]),   .b4(a[4] & b[12]),   .b5(a[5] & b[12]),   .b6(a[6] & b[12]),   .b7(a[7] & b[12]),
			        .b8(a[8] & b[12]),   .b9(a[9] & b[12]),   .b10(a[10] & b[12]), .b11(a[12] & b[12]), .b12(a[12] & b[12]), .b13(a[13] & b[12]), .b14(a[14] & b[12]), .b15(a[15] & b[12]),
			        .b16(a[16] & b[12]), .b17(a[17] & b[12]), .b18(a[18] & b[12]), .b19(a[19] & b[12]), .b20(a[20] & b[12]), .b21(a[21] & b[12]), .b22(a[22] & b[12]), .b23(a[23] & b[12]),
	                        .b24(a[24] & b[12]), .b25(a[25] & b[12]), .b26(a[26] & b[12]), .b27(a[27] & b[12]), .b28(a[28] & b[12]), .b29(a[29] & b[12]), .b30(a[30] & b[12]), .b31(a[31] & b[12]),	  
	          .cin(1'b0), .cout(carry12));

fullAdder32b fa13 (.sum(sum13), .a0(sum12[1]),   .a1(sum12[2]),   .a2(sum12[3]),   .a3(sum12[4]),   .a4(sum12[5]),   .a5(sum12[6]),   .a6(sum12[7]),   .a7(sum12[8]),   .a8(sum12[9]),   .a9(sum12[10]),  .a10(sum12[11]), 
		                .a11(sum12[12]), .a12(sum12[13]), .a13(sum12[14]), .a14(sum12[15]), .a15(sum12[16]), .a16(sum12[17]), .a17(sum12[18]), .a18(sum12[19]), .a19(sum12[20]), .a20(sum12[21]), .a21(sum12[22]),
			        .a22(sum12[23]), .a23(sum12[24]), .a24(sum12[25]), .a25(sum12[26]), .a26(sum12[27]), .a27(sum12[28]), .a28(sum12[29]), .a29(sum12[30]), .a30(sum12[31]), .a31(carry12),

			        .b0(a[0] & b[13]),   .b1(a[1] & b[13]),   .b2(a[2] & b[13]),   .b3(a[3] & b[13]),   .b4(a[4] & b[13]),   .b5(a[5] & b[13]),   .b6(a[6] & b[13]),   .b7(a[7] & b[13]),
			        .b8(a[8] & b[13]),   .b9(a[9] & b[13]),   .b10(a[10] & b[13]), .b11(a[12] & b[13]), .b12(a[12] & b[13]), .b13(a[13] & b[13]), .b14(a[14] & b[13]), .b15(a[15] & b[13]),
			        .b16(a[16] & b[13]), .b17(a[17] & b[13]), .b18(a[18] & b[13]), .b19(a[19] & b[13]), .b20(a[20] & b[13]), .b21(a[21] & b[13]), .b22(a[22] & b[13]), .b23(a[23] & b[13]),
	                        .b24(a[24] & b[13]), .b25(a[25] & b[13]), .b26(a[26] & b[13]), .b27(a[27] & b[13]), .b28(a[28] & b[13]), .b29(a[29] & b[13]), .b30(a[30] & b[13]), .b31(a[31] & b[13]),	  
	          .cin(1'b0), .cout(carry13));

fullAdder32b fa14 (.sum(sum14), .a0(sum13[1]),   .a1(sum13[2]),   .a2(sum13[3]),   .a3(sum13[4]),   .a4(sum13[5]),   .a5(sum13[6]),   .a6(sum13[7]),   .a7(sum13[8]),   .a8(sum13[9]),   .a9(sum13[10]),  .a10(sum13[11]), 
		                .a11(sum13[12]), .a12(sum13[13]), .a13(sum13[14]), .a14(sum13[15]), .a15(sum13[16]), .a16(sum13[17]), .a17(sum13[18]), .a18(sum13[19]), .a19(sum13[20]), .a20(sum13[21]), .a21(sum13[22]),
			        .a22(sum13[23]), .a23(sum13[24]), .a24(sum13[25]), .a25(sum13[26]), .a26(sum13[27]), .a27(sum13[28]), .a28(sum13[29]), .a29(sum13[30]), .a30(sum13[31]), .a31(carry13), 

			        .b0(a[0] & b[14]),   .b1(a[1] & b[14]),   .b2(a[2] & b[14]),   .b3(a[3] & b[14]),   .b4(a[4] & b[14]),   .b5(a[5] & b[14]),   .b6(a[6] & b[14]),   .b7(a[7] & b[14]),
			        .b8(a[8] & b[14]),   .b9(a[9] & b[14]),   .b10(a[10] & b[14]), .b11(a[12] & b[14]), .b12(a[12] & b[14]), .b13(a[13] & b[14]), .b14(a[14] & b[14]), .b15(a[15] & b[14]),
			        .b16(a[16] & b[14]), .b17(a[17] & b[14]), .b18(a[18] & b[14]), .b19(a[19] & b[14]), .b20(a[20] & b[14]), .b21(a[21] & b[14]), .b22(a[22] & b[14]), .b23(a[23] & b[14]),
	                        .b24(a[24] & b[14]), .b25(a[25] & b[14]), .b26(a[26] & b[14]), .b27(a[27] & b[14]), .b28(a[28] & b[14]), .b29(a[29] & b[14]), .b30(a[30] & b[14]), .b31(a[31] & b[14]),	  
	          .cin(1'b0), .cout(carry14));

fullAdder32b fa15 (.sum(sum15), .a0(sum14[1]),   .a1(sum14[2]),   .a2(sum14[3]),   .a3(sum14[4]),   .a4(sum14[5]),   .a5(sum14[6]),   .a6(sum14[7]),   .a7(sum14[8]),   .a8(sum14[9]),   .a9(sum14[10]),  .a10(sum14[11]), 
		                .a11(sum14[12]), .a12(sum14[13]), .a13(sum14[14]), .a14(sum14[15]), .a15(sum14[16]), .a16(sum14[17]), .a17(sum14[18]), .a18(sum14[19]), .a19(sum14[20]), .a20(sum14[21]), .a21(sum14[22]),
			        .a22(sum14[23]), .a23(sum14[24]), .a24(sum14[25]), .a25(sum14[26]), .a26(sum14[27]), .a27(sum14[28]), .a28(sum14[29]), .a29(sum14[30]), .a30(sum14[31]), .a31(carry14), 

			        .b0(a[0] & b[15]),   .b1(a[1] & b[15]),   .b2(a[2] & b[15]),   .b3(a[3] & b[15]),   .b4(a[4] & b[15]),   .b5(a[5] & b[15]),   .b6(a[6] & b[15]),   .b7(a[7] & b[15]),
			        .b8(a[8] & b[15]),   .b9(a[9] & b[15]),   .b10(a[10] & b[15]), .b11(a[12] & b[15]), .b12(a[12] & b[15]), .b13(a[13] & b[15]), .b14(a[14] & b[15]), .b15(a[15] & b[15]),
			        .b16(a[16] & b[15]), .b17(a[17] & b[15]), .b18(a[18] & b[15]), .b19(a[19] & b[15]), .b20(a[20] & b[15]), .b21(a[21] & b[15]), .b22(a[22] & b[15]), .b23(a[23] & b[15]),
	                        .b24(a[24] & b[15]), .b25(a[25] & b[15]), .b26(a[26] & b[15]), .b27(a[27] & b[15]), .b28(a[28] & b[15]), .b29(a[29] & b[15]), .b30(a[30] & b[15]), .b31(a[31] & b[15]),	  
	          .cin(1'b0), .cout(carry15));

fullAdder32b fa16 (.sum(sum16), .a0(sum15[1]),   .a1(sum15[2]),   .a2(sum15[3]),   .a3(sum15[4]),   .a4(sum15[5]),   .a5(sum15[6]),   .a6(sum15[7]),   .a7(sum15[8]),   .a8(sum15[9]),   .a9(sum15[10]),  .a10(sum15[11]), 
		                .a11(sum15[12]), .a12(sum15[13]), .a13(sum15[14]), .a14(sum15[15]), .a15(sum15[16]), .a16(sum15[17]), .a17(sum15[18]), .a18(sum15[19]), .a19(sum15[20]), .a20(sum15[21]), .a21(sum15[22]),
			        .a22(sum15[23]), .a23(sum15[24]), .a24(sum15[25]), .a25(sum15[26]), .a26(sum15[27]), .a27(sum15[28]), .a28(sum15[29]), .a29(sum15[30]), .a30(sum15[31]), .a31(carry15), 

			        .b0(a[0] & b[16]),   .b1(a[1] & b[16]),   .b2(a[2] & b[16]),   .b3(a[3] & b[16]),   .b4(a[4] & b[16]),   .b5(a[5] & b[16]),   .b6(a[6] & b[16]),   .b7(a[7] & b[16]),
			        .b8(a[8] & b[16]),   .b9(a[9] & b[16]),   .b10(a[10] & b[16]), .b11(a[12] & b[16]), .b12(a[12] & b[16]), .b13(a[13] & b[16]), .b14(a[14] & b[16]), .b15(a[15] & b[16]),
			        .b16(a[16] & b[16]), .b17(a[17] & b[16]), .b18(a[18] & b[16]), .b19(a[19] & b[16]), .b20(a[20] & b[16]), .b21(a[21] & b[16]), .b22(a[22] & b[16]), .b23(a[23] & b[16]),
	                        .b24(a[24] & b[16]), .b25(a[25] & b[16]), .b26(a[26] & b[16]), .b27(a[27] & b[16]), .b28(a[28] & b[16]), .b29(a[29] & b[16]), .b30(a[30] & b[16]), .b31(a[31] & b[16]),	  
	          .cin(1'b0), .cout(carry16));

fullAdder32b fa17 (.sum(sum17), .a0(sum16[1]),   .a1(sum16[2]),   .a2(sum16[3]),   .a3(sum16[4]),   .a4(sum16[5]),   .a5(sum16[6]),   .a6(sum16[7]),   .a7(sum16[8]),   .a8(sum16[9]),   .a9(sum16[10]),  .a10(sum16[11]), 
		                .a11(sum16[12]), .a12(sum16[13]), .a13(sum16[14]), .a14(sum16[15]), .a15(sum16[16]), .a16(sum16[17]), .a17(sum16[18]), .a18(sum16[19]), .a19(sum16[20]), .a20(sum16[21]), .a21(sum16[22]),
			        .a22(sum16[23]), .a23(sum16[24]), .a24(sum16[25]), .a25(sum16[26]), .a26(sum16[27]), .a27(sum16[28]), .a28(sum16[29]), .a29(sum16[30]), .a30(sum16[31]), .a31(carry16), 

			        .b0(a[0] & b[17]),   .b1(a[1] & b[17]),   .b2(a[2] & b[17]),   .b3(a[3] & b[17]),   .b4(a[4] & b[17]),   .b5(a[5] & b[17]),   .b6(a[6] & b[17]),   .b7(a[7] & b[17]),
			        .b8(a[8] & b[17]),   .b9(a[9] & b[17]),   .b10(a[10] & b[17]), .b11(a[12] & b[17]), .b12(a[12] & b[17]), .b13(a[13] & b[17]), .b14(a[14] & b[17]), .b15(a[15] & b[17]),
			        .b16(a[16] & b[17]), .b17(a[17] & b[17]), .b18(a[18] & b[17]), .b19(a[19] & b[17]), .b20(a[20] & b[17]), .b21(a[21] & b[17]), .b22(a[22] & b[17]), .b23(a[23] & b[17]),
	                        .b24(a[24] & b[17]), .b25(a[25] & b[17]), .b26(a[26] & b[17]), .b27(a[27] & b[17]), .b28(a[28] & b[17]), .b29(a[29] & b[17]), .b30(a[30] & b[17]), .b31(a[31] & b[17]),	  
	          .cin(1'b0), .cout(carry17));

fullAdder32b fa18 (.sum(sum18), .a0(sum17[1]),   .a1(sum17[2]),   .a2(sum17[3]),   .a3(sum17[4]),   .a4(sum17[5]),   .a5(sum17[6]),   .a6(sum17[7]),   .a7(sum17[8]),   .a8(sum17[9]),   .a9(sum17[10]),  .a10(sum17[11]), 
		                .a11(sum17[12]), .a12(sum17[13]), .a13(sum17[14]), .a14(sum17[15]), .a15(sum17[16]), .a16(sum17[17]), .a17(sum17[18]), .a18(sum17[19]), .a19(sum17[20]), .a20(sum17[21]), .a21(sum17[22]),
			        .a22(sum17[23]), .a23(sum17[24]), .a24(sum17[25]), .a25(sum17[26]), .a26(sum17[27]), .a27(sum17[28]), .a28(sum17[29]), .a29(sum17[30]), .a30(sum17[31]), .a31(carry17), 

			        .b0(a[0] & b[18]),   .b1(a[1] & b[18]),   .b2(a[2] & b[18]),   .b3(a[3] & b[18]),   .b4(a[4] & b[18]),   .b5(a[5] & b[18]),   .b6(a[6] & b[18]),   .b7(a[7] & b[18]),
			        .b8(a[8] & b[18]),   .b9(a[9] & b[18]),   .b10(a[10] & b[18]), .b11(a[12] & b[18]), .b12(a[12] & b[18]), .b13(a[13] & b[18]), .b14(a[14] & b[18]), .b15(a[15] & b[18]),
			        .b16(a[16] & b[18]), .b17(a[17] & b[18]), .b18(a[18] & b[18]), .b19(a[19] & b[18]), .b20(a[20] & b[18]), .b21(a[21] & b[18]), .b22(a[22] & b[18]), .b23(a[23] & b[18]),
	                        .b24(a[24] & b[18]), .b25(a[25] & b[18]), .b26(a[26] & b[18]), .b27(a[27] & b[18]), .b28(a[28] & b[18]), .b29(a[29] & b[18]), .b30(a[30] & b[18]), .b31(a[31] & b[18]),	  
	          .cin(1'b0), .cout(carry18));

fullAdder32b fa19 (.sum(sum19), .a0(sum18[1]),   .a1(sum18[2]),   .a2(sum18[3]),   .a3(sum18[4]),   .a4(sum18[5]),   .a5(sum18[6]),   .a6(sum18[7]),   .a7(sum18[8]),   .a8(sum18[9]),   .a9(sum18[10]),  .a10(sum18[11]), 
		                .a11(sum18[12]), .a12(sum18[13]), .a13(sum18[14]), .a14(sum18[15]), .a15(sum18[16]), .a16(sum18[17]), .a17(sum18[18]), .a18(sum18[19]), .a19(sum18[20]), .a20(sum18[21]), .a21(sum18[22]),
			        .a22(sum18[23]), .a23(sum18[24]), .a24(sum18[25]), .a25(sum18[26]), .a26(sum18[27]), .a27(sum18[28]), .a28(sum18[29]), .a29(sum18[30]), .a30(sum18[31]), .a31(carry18), 

			        .b0(a[0] & b[19]),   .b1(a[1] & b[19]),   .b2(a[2] & b[19]),   .b3(a[3] & b[19]),   .b4(a[4] & b[11]),   .b5(a[5] & b[19]),   .b6(a[6] & b[19]),   .b7(a[7] & b[19]),
			        .b8(a[8] & b[19]),   .b9(a[9] & b[19]),   .b10(a[10] & b[19]), .b11(a[12] & b[19]), .b12(a[12] & b[19]), .b13(a[13] & b[19]), .b14(a[14] & b[19]), .b15(a[15] & b[19]),
			        .b16(a[16] & b[19]), .b17(a[17] & b[19]), .b18(a[18] & b[19]), .b19(a[19] & b[19]), .b20(a[20] & b[19]), .b21(a[21] & b[19]), .b22(a[22] & b[19]), .b23(a[23] & b[19]),
	                        .b24(a[24] & b[19]), .b25(a[25] & b[19]), .b26(a[26] & b[19]), .b27(a[27] & b[19]), .b28(a[28] & b[19]), .b29(a[29] & b[19]), .b30(a[30] & b[19]), .b31(a[31] & b[19]),	  
	          .cin(1'b0), .cout(carry19));

fullAdder32b fa20 (.sum(sum20), .a0(sum19[1]),   .a1(sum19[2]),   .a2(sum19[3]),   .a3(sum19[4]),   .a4(sum19[5]),   .a5(sum19[6]),   .a6(sum19[7]),   .a7(sum19[8]),   .a8(sum19[9]),   .a9(sum19[10]),  .a10(sum19[11]), 
		                .a11(sum19[12]), .a12(sum19[13]), .a13(sum19[14]), .a14(sum19[15]), .a15(sum19[16]), .a16(sum19[17]), .a17(sum19[18]), .a18(sum19[19]), .a19(sum19[20]), .a20(sum19[21]), .a21(sum19[22]),
			        .a22(sum19[23]), .a23(sum19[24]), .a24(sum19[25]), .a25(sum19[26]), .a26(sum19[27]), .a27(sum19[28]), .a28(sum19[29]), .a29(sum19[30]), .a30(sum19[31]), .a31(carry19), 

			        .b0(a[0] & b[20]),   .b1(a[1] & b[20]),   .b2(a[2] & b[20]),   .b3(a[3] & b[20]),   .b4(a[4] & b[20]),   .b5(a[5] & b[20]),   .b6(a[6] & b[20]),   .b7(a[7] & b[20]),
			        .b8(a[8] & b[20]),   .b9(a[9] & b[20]),   .b10(a[10] & b[20]), .b11(a[12] & b[20]), .b12(a[12] & b[20]), .b13(a[13] & b[20]), .b14(a[14] & b[20]), .b15(a[15] & b[20]),
			        .b16(a[16] & b[20]), .b17(a[17] & b[20]), .b18(a[18] & b[20]), .b19(a[19] & b[20]), .b20(a[20] & b[20]), .b21(a[21] & b[20]), .b22(a[22] & b[20]), .b23(a[23] & b[20]),
	                        .b24(a[24] & b[20]), .b25(a[25] & b[20]), .b26(a[26] & b[20]), .b27(a[27] & b[20]), .b28(a[28] & b[20]), .b29(a[29] & b[20]), .b30(a[30] & b[20]), .b31(a[31] & b[20]),	  
	          .cin(1'b0), .cout(carry20));


fullAdder32b fa21 (.sum(sum21), .a0(sum20[1]),   .a1(sum20[2]),   .a2(sum20[3]),   .a3(sum20[4]),   .a4(sum20[5]),   .a5(sum20[6]),   .a6(sum20[7]),   .a7(sum20[8]),   .a8(sum20[9]),   .a9(sum20[10]),  .a10(sum20[11]), 
		                .a11(sum20[12]), .a12(sum20[13]), .a13(sum20[14]), .a14(sum20[15]), .a15(sum20[16]), .a16(sum20[17]), .a17(sum20[18]), .a18(sum20[19]), .a19(sum20[20]), .a20(sum20[21]), .a21(sum20[22]),
			        .a22(sum20[23]), .a23(sum20[24]), .a24(sum20[25]), .a25(sum20[26]), .a26(sum20[27]), .a27(sum20[28]), .a28(sum20[29]), .a29(sum20[30]), .a30(sum20[31]), .a31(carry20), 

			        .b0(a[0] & b[21]),   .b1(a[1] & b[21]),   .b2(a[2] & b[21]),   .b3(a[3] & b[21]),   .b4(a[4] & b[21]),   .b5(a[5] & b[21]),   .b6(a[6] & b[21]),   .b7(a[7] & b[21]),
			        .b8(a[8] & b[21]),   .b9(a[9] & b[21]),   .b10(a[10] & b[21]), .b11(a[12] & b[21]), .b12(a[12] & b[21]), .b13(a[13] & b[21]), .b14(a[14] & b[21]), .b15(a[15] & b[21]),
			        .b16(a[16] & b[21]), .b17(a[17] & b[21]), .b18(a[18] & b[21]), .b19(a[19] & b[21]), .b20(a[20] & b[21]), .b21(a[21] & b[21]), .b22(a[22] & b[21]), .b23(a[23] & b[21]),
	                        .b24(a[24] & b[21]), .b25(a[25] & b[21]), .b26(a[26] & b[21]), .b27(a[27] & b[21]), .b28(a[28] & b[21]), .b29(a[29] & b[21]), .b30(a[30] & b[21]), .b31(a[31] & b[21]),	  
	          .cin(1'b0), .cout(carry21));

fullAdder32b fa22 (.sum(sum22), .a0(sum21[1]),   .a1(sum21[2]),   .a2(sum21[3]),   .a3(sum21[4]),   .a4(sum21[5]),   .a5(sum21[6]),   .a6(sum21[7]),   .a7(sum21[8]),   .a8(sum21[9]),   .a9(sum21[10]),  .a10(sum21[11]), 
		                .a11(sum21[12]), .a12(sum21[13]), .a13(sum21[14]), .a14(sum21[15]), .a15(sum21[16]), .a16(sum21[17]), .a17(sum21[18]), .a18(sum21[19]), .a19(sum21[20]), .a20(sum21[21]), .a21(sum21[22]),
			        .a22(sum21[23]), .a23(sum21[24]), .a24(sum21[25]), .a25(sum21[26]), .a26(sum21[27]), .a27(sum21[28]), .a28(sum21[29]), .a29(sum21[30]), .a30(sum21[31]), .a31(carry21), 

			        .b0(a[0] & b[22]),   .b1(a[1] & b[22]),   .b2(a[2] & b[22]),   .b3(a[3] & b[22]),   .b4(a[4] & b[22]),   .b5(a[5] & b[22]),   .b6(a[6] & b[22]),   .b7(a[7] & b[22]),
			        .b8(a[8] & b[22]),   .b9(a[9] & b[22]),   .b10(a[10] & b[22]), .b11(a[12] & b[22]), .b12(a[12] & b[22]), .b13(a[13] & b[22]), .b14(a[14] & b[22]), .b15(a[15] & b[22]),
			        .b16(a[16] & b[22]), .b17(a[17] & b[22]), .b18(a[18] & b[22]), .b19(a[19] & b[22]), .b20(a[20] & b[22]), .b21(a[21] & b[22]), .b22(a[22] & b[22]), .b23(a[23] & b[22]),
	                        .b24(a[24] & b[22]), .b25(a[25] & b[22]), .b26(a[26] & b[22]), .b27(a[27] & b[22]), .b28(a[28] & b[22]), .b29(a[29] & b[22]), .b30(a[30] & b[22]), .b31(a[31] & b[22]),	  
	          .cin(1'b0), .cout(carry22));
	  
fullAdder32b fa23 (.sum(sum23), .a0(sum22[1]),   .a1(sum22[2]),   .a2(sum22[3]),   .a3(sum22[4]),   .a4(sum22[5]),   .a5(sum22[6]),   .a6(sum22[7]),   .a7(sum22[8]),   .a8(sum22[9]),   .a9(sum22[10]),  .a10(sum22[11]), 
		                .a11(sum22[12]), .a12(sum22[13]), .a13(sum22[14]), .a14(sum22[15]), .a15(sum22[16]), .a16(sum22[17]), .a17(sum22[18]), .a18(sum22[19]), .a19(sum22[20]), .a20(sum22[21]), .a21(sum22[22]),
			        .a22(sum22[23]), .a23(sum22[24]), .a24(sum22[25]), .a25(sum22[26]), .a26(sum22[27]), .a27(sum22[28]), .a28(sum22[29]), .a29(sum22[30]), .a30(sum22[31]), .a31(carry22), 

			        .b0(a[0] & b[23]),   .b1(a[1] & b[23]),   .b2(a[2] & b[23]),   .b3(a[3] & b[23]),   .b4(a[4] & b[23]),   .b5(a[5] & b[23]),   .b6(a[6] & b[23]),   .b7(a[7] & b[23]),
			        .b8(a[8] & b[23]),   .b9(a[9] & b[23]),   .b10(a[10] & b[23]), .b11(a[12] & b[23]), .b12(a[12] & b[23]), .b13(a[13] & b[23]), .b14(a[14] & b[23]), .b15(a[15] & b[23]),
			        .b16(a[16] & b[23]), .b17(a[17] & b[23]), .b18(a[18] & b[23]), .b19(a[19] & b[23]), .b20(a[20] & b[23]), .b21(a[21] & b[23]), .b22(a[22] & b[23]), .b23(a[23] & b[23]),
	                        .b24(a[24] & b[23]), .b25(a[25] & b[23]), .b26(a[26] & b[23]), .b27(a[27] & b[23]), .b28(a[28] & b[23]), .b29(a[29] & b[23]), .b30(a[30] & b[23]), .b31(a[31] & b[23]),	  
	          .cin(1'b0), .cout(carry23));
	  
fullAdder32b fa24 (.sum(sum24), .a0(sum23[1]),   .a1(sum23[2]),   .a2(sum23[3]),   .a3(sum23[4]),   .a4(sum23[5]),   .a5(sum23[6]),   .a6(sum23[7]),   .a7(sum23[8]),   .a8(sum23[9]),   .a9(sum23[10]),  .a10(sum23[11]), 
		                .a11(sum23[12]), .a12(sum23[13]), .a13(sum23[14]), .a14(sum23[15]), .a15(sum23[16]), .a16(sum23[17]), .a17(sum23[18]), .a18(sum23[19]), .a19(sum23[20]), .a20(sum23[21]), .a21(sum23[22]),
			        .a22(sum23[23]), .a23(sum23[24]), .a24(sum23[25]), .a25(sum23[26]), .a26(sum23[27]), .a27(sum23[28]), .a28(sum23[29]), .a29(sum23[30]), .a30(sum23[31]), .a31(carry23), 

			        .b0(a[0] & b[24]),   .b1(a[1] & b[24]),   .b2(a[2] & b[24]),   .b3(a[3] & b[24]),   .b4(a[4] & b[24]),   .b5(a[5] & b[24]),   .b6(a[6] & b[24]),   .b7(a[7] & b[24]),
			        .b8(a[8] & b[24]),   .b9(a[9] & b[24]),   .b10(a[10] & b[24]), .b11(a[12] & b[24]), .b12(a[12] & b[24]), .b13(a[13] & b[24]), .b14(a[14] & b[24]), .b15(a[15] & b[24]),
			        .b16(a[16] & b[24]), .b17(a[17] & b[24]), .b18(a[18] & b[24]), .b19(a[19] & b[24]), .b20(a[20] & b[24]), .b21(a[21] & b[24]), .b22(a[22] & b[24]), .b23(a[23] & b[24]),
	                        .b24(a[24] & b[24]), .b25(a[25] & b[24]), .b26(a[26] & b[24]), .b27(a[27] & b[24]), .b28(a[28] & b[24]), .b29(a[29] & b[24]), .b30(a[30] & b[24]), .b31(a[31] & b[24]),	  
	          .cin(1'b0), .cout(carry24));


fullAdder32b fa25 (.sum(sum25), .a0(sum24[1]),   .a1(sum24[2]),   .a2(sum24[3]),   .a3(sum24[4]),   .a4(sum24[5]),   .a5(sum24[6]),   .a6(sum24[7]),   .a7(sum24[8]),   .a8(sum24[9]),   .a9(sum24[10]),  .a10(sum24[11]), 
		                .a11(sum24[12]), .a12(sum24[13]), .a13(sum24[14]), .a14(sum24[15]), .a15(sum24[16]), .a16(sum24[17]), .a17(sum24[18]), .a18(sum24[19]), .a19(sum24[20]), .a20(sum24[21]), .a21(sum24[22]),
			        .a22(sum24[23]), .a23(sum24[24]), .a24(sum24[25]), .a25(sum24[26]), .a26(sum24[27]), .a27(sum24[28]), .a28(sum24[29]), .a29(sum24[30]), .a30(sum24[31]), .a31(carry24), 

			        .b0(a[0] & b[25]),   .b1(a[1] & b[25]),   .b2(a[2] & b[25]),   .b3(a[3] & b[25]),   .b4(a[4] & b[25]),   .b5(a[5] & b[25]),   .b6(a[6] & b[25]),   .b7(a[7] & b[25]),
			        .b8(a[8] & b[25]),   .b9(a[9] & b[25]),   .b10(a[10] & b[25]), .b11(a[12] & b[25]), .b12(a[12] & b[25]), .b13(a[13] & b[25]), .b14(a[14] & b[25]), .b15(a[15] & b[25]),
			        .b16(a[16] & b[25]), .b17(a[17] & b[25]), .b18(a[18] & b[25]), .b19(a[19] & b[25]), .b20(a[20] & b[25]), .b21(a[21] & b[25]), .b22(a[22] & b[25]), .b23(a[23] & b[25]),
	                        .b24(a[24] & b[25]), .b25(a[25] & b[25]), .b26(a[26] & b[25]), .b27(a[27] & b[25]), .b28(a[28] & b[25]), .b29(a[29] & b[25]), .b30(a[30] & b[25]), .b31(a[31] & b[25]),	  
	          .cin(1'b0), .cout(carry25));
	  	  
fullAdder32b fa26 (.sum(sum26), .a0(sum25[1]),   .a1(sum25[2]),   .a2(sum25[3]),   .a3(sum25[4]),   .a4(sum25[5]),   .a5(sum25[6]),   .a6(sum25[7]),   .a7(sum25[8]),   .a8(sum25[9]),   .a9(sum25[10]),  .a10(sum25[11]), 
		                .a11(sum25[12]), .a12(sum25[13]), .a13(sum25[14]), .a14(sum25[15]), .a15(sum25[16]), .a16(sum25[17]), .a17(sum25[18]), .a18(sum25[19]), .a19(sum25[20]), .a20(sum25[21]), .a21(sum25[22]),
			        .a22(sum25[23]), .a23(sum25[24]), .a24(sum25[25]), .a25(sum25[26]), .a26(sum25[27]), .a27(sum25[28]), .a28(sum25[29]), .a29(sum25[30]), .a30(sum25[31]), .a31(carry25), 

			        .b0(a[0] & b[26]),   .b1(a[1] & b[26]),   .b2(a[2] & b[26]),   .b3(a[3] & b[26]),   .b4(a[4] & b[26]),   .b5(a[5] & b[26]),   .b6(a[6] & b[26]),   .b7(a[7] & b[26]),
			        .b8(a[8] & b[26]),   .b9(a[9] & b[26]),   .b10(a[10] & b[26]), .b11(a[12] & b[26]), .b12(a[12] & b[26]), .b13(a[13] & b[26]), .b14(a[14] & b[26]), .b15(a[15] & b[26]),
			        .b16(a[16] & b[26]), .b17(a[17] & b[26]), .b18(a[18] & b[26]), .b19(a[19] & b[26]), .b20(a[20] & b[26]), .b21(a[21] & b[26]), .b22(a[22] & b[26]), .b23(a[23] & b[26]),
	                        .b24(a[24] & b[26]), .b25(a[25] & b[26]), .b26(a[26] & b[26]), .b27(a[27] & b[26]), .b28(a[28] & b[26]), .b29(a[29] & b[26]), .b30(a[30] & b[26]), .b31(a[31] & b[26]),	  
	          .cin(1'b0), .cout(carry26));

fullAdder32b fa27 (.sum(sum27), .a0(sum26[1]),   .a1(sum26[2]),   .a2(sum26[3]),   .a3(sum26[4]),   .a4(sum26[5]),   .a5(sum26[6]),   .a6(sum26[7]),   .a7(sum26[8]),   .a8(sum26[9]),   .a9(sum26[10]),  .a10(sum26[11]), 
		                .a11(sum26[12]), .a12(sum26[13]), .a13(sum26[14]), .a14(sum26[15]), .a15(sum26[16]), .a16(sum26[17]), .a17(sum26[18]), .a18(sum26[19]), .a19(sum26[20]), .a20(sum26[21]), .a21(sum26[22]),
			        .a22(sum26[23]), .a23(sum26[24]), .a24(sum26[25]), .a25(sum26[26]), .a26(sum26[27]), .a27(sum26[28]), .a28(sum26[29]), .a29(sum26[30]), .a30(sum26[31]), .a31(carry26), 

			        .b0(a[0] & b[27]),   .b1(a[1] & b[27]),   .b2(a[2] & b[27]),   .b3(a[3] & b[27]),   .b4(a[4] & b[27]),   .b5(a[5] & b[27]),   .b6(a[6] & b[27]),   .b7(a[7] & b[27]),
			        .b8(a[8] & b[27]),   .b9(a[9] & b[27]),   .b10(a[10] & b[27]), .b11(a[12] & b[27]), .b12(a[12] & b[27]), .b13(a[13] & b[27]), .b14(a[14] & b[27]), .b15(a[15] & b[27]),
			        .b16(a[16] & b[27]), .b17(a[17] & b[27]), .b18(a[18] & b[27]), .b19(a[19] & b[27]), .b20(a[20] & b[27]), .b21(a[21] & b[27]), .b22(a[22] & b[27]), .b23(a[23] & b[27]),
	                        .b24(a[24] & b[27]), .b25(a[25] & b[27]), .b26(a[26] & b[27]), .b27(a[27] & b[27]), .b28(a[28] & b[27]), .b29(a[29] & b[27]), .b30(a[30] & b[27]), .b31(a[31] & b[27]),	  
	          .cin(1'b0), .cout(carry27));

fullAdder32b fa28 (.sum(sum28), .a0(sum27[1]),   .a1(sum27[2]),   .a2(sum27[3]),   .a3(sum27[4]),   .a4(sum27[5]),   .a5(sum27[6]),   .a6(sum27[7]),   .a7(sum27[8]),   .a8(sum27[9]),   .a9(sum27[10]),  .a10(sum27[11]), 
		                .a11(sum27[12]), .a12(sum27[13]), .a13(sum27[14]), .a14(sum27[15]), .a15(sum27[16]), .a16(sum27[17]), .a17(sum27[18]), .a18(sum27[19]), .a19(sum27[20]), .a20(sum27[21]), .a21(sum27[22]),
			        .a22(sum27[23]), .a23(sum27[24]), .a24(sum27[25]), .a25(sum27[26]), .a26(sum27[27]), .a27(sum27[28]), .a28(sum27[29]), .a29(sum27[30]), .a30(sum27[31]), .a31(carry27), 

			        .b0(a[0] & b[28]),   .b1(a[1] & b[28]),   .b2(a[2] & b[28]),   .b3(a[3] & b[28]),   .b4(a[4] & b[28]),   .b5(a[5] & b[28]),   .b6(a[6] & b[28]),   .b7(a[7] & b[28]),
			        .b8(a[8] & b[28]),   .b9(a[9] & b[28]),   .b10(a[10] & b[28]), .b11(a[12] & b[28]), .b12(a[12] & b[28]), .b13(a[13] & b[28]), .b14(a[14] & b[28]), .b15(a[15] & b[28]),
			        .b16(a[16] & b[28]), .b17(a[17] & b[28]), .b18(a[18] & b[28]), .b19(a[19] & b[28]), .b20(a[20] & b[28]), .b21(a[21] & b[28]), .b22(a[22] & b[28]), .b23(a[23] & b[28]),
	                        .b24(a[24] & b[28]), .b25(a[25] & b[28]), .b26(a[26] & b[28]), .b27(a[27] & b[28]), .b28(a[28] & b[28]), .b29(a[29] & b[28]), .b30(a[30] & b[28]), .b31(a[31] & b[28]),	  
	          .cin(1'b0), .cout(carry28));


fullAdder32b fa29 (.sum(sum29), .a0(sum28[1]),   .a1(sum28[2]),   .a2(sum28[3]),   .a3(sum28[4]),   .a4(sum28[5]),   .a5(sum28[6]),   .a6(sum28[7]),   .a7(sum28[8]),   .a8(sum28[9]),   .a9(sum28[10]),  .a10(sum28[11]), 
		                .a11(sum28[12]), .a12(sum28[13]), .a13(sum28[14]), .a14(sum28[15]), .a15(sum28[16]), .a16(sum28[17]), .a17(sum28[18]), .a18(sum28[19]), .a19(sum28[20]), .a20(sum28[21]), .a21(sum28[22]),
			        .a22(sum28[23]), .a23(sum28[24]), .a24(sum28[25]), .a25(sum28[26]), .a26(sum28[27]), .a27(sum28[28]), .a28(sum28[29]), .a29(sum28[30]), .a30(sum28[31]), .a31(carry28), 

			        .b0(a[0] & b[29]),   .b1(a[1] & b[29]),   .b2(a[2] & b[29]),   .b3(a[3] & b[29]),   .b4(a[4] & b[29]),   .b5(a[5] & b[29]),   .b6(a[6] & b[29]),   .b7(a[7] & b[29]),
			        .b8(a[8] & b[29]),   .b9(a[9] & b[29]),   .b10(a[10] & b[29]), .b11(a[12] & b[29]), .b12(a[12] & b[29]), .b13(a[13] & b[29]), .b14(a[14] & b[29]), .b15(a[15] & b[29]),
			        .b16(a[16] & b[29]), .b17(a[17] & b[29]), .b18(a[18] & b[29]), .b19(a[19] & b[29]), .b20(a[20] & b[29]), .b21(a[21] & b[29]), .b22(a[22] & b[29]), .b23(a[23] & b[29]),
	                        .b24(a[24] & b[29]), .b25(a[25] & b[29]), .b26(a[26] & b[29]), .b27(a[27] & b[29]), .b28(a[28] & b[29]), .b29(a[29] & b[29]), .b30(a[30] & b[29]), .b31(a[31] & b[29]),	  
	          .cin(1'b0), .cout(carry29));

fullAdder32b fa30 (.sum(sum30), .a0(sum29[1]),   .a1(sum29[2]),   .a2(sum29[3]),   .a3(sum29[4]),   .a4(sum29[5]),   .a5(sum29[6]),   .a6(sum29[7]),   .a7(sum29[8]),   .a8(sum29[9]),   .a9(sum29[10]),  .a10(sum29[11]), 
		                .a11(sum29[12]), .a12(sum29[13]), .a13(sum29[14]), .a14(sum29[15]), .a15(sum29[16]), .a16(sum29[17]), .a17(sum29[18]), .a18(sum29[19]), .a19(sum29[20]), .a20(sum29[21]), .a21(sum29[22]),
			        .a22(sum29[23]), .a23(sum29[24]), .a24(sum29[25]), .a25(sum29[26]), .a26(sum29[27]), .a27(sum29[28]), .a28(sum29[29]), .a29(sum29[30]), .a30(sum29[31]), .a31(carry29), 

			        .b0(a[0] & b[30]),   .b1(a[1] & b[30]),   .b2(a[2] & b[30]),   .b3(a[3] & b[30]),   .b4(a[4] & b[30]),   .b5(a[5] & b[30]),   .b6(a[6] & b[30]),   .b7(a[7] & b[30]),
			        .b8(a[8] & b[30]),   .b9(a[9] & b[30]),   .b10(a[10] & b[30]), .b11(a[12] & b[30]), .b12(a[12] & b[30]), .b13(a[13] & b[30]), .b14(a[14] & b[30]), .b15(a[15] & b[30]),
			        .b16(a[16] & b[30]), .b17(a[17] & b[30]), .b18(a[18] & b[30]), .b19(a[19] & b[30]), .b20(a[20] & b[30]), .b21(a[21] & b[30]), .b22(a[22] & b[30]), .b23(a[23] & b[30]),
	                        .b24(a[24] & b[30]), .b25(a[25] & b[30]), .b26(a[26] & b[30]), .b27(a[27] & b[30]), .b28(a[28] & b[30]), .b29(a[29] & b[30]), .b30(a[30] & b[30]), .b31(a[31] & b[30]),	  
	          .cin(1'b0), .cout(carry30));

fullAdder32b fa31 (.sum(sum31), .a0(sum30[1]),   .a1(sum30[2]),   .a2(sum30[3]),   .a3(sum30[4]),   .a4(sum30[5]),   .a5(sum30[6]),   .a6(sum30[7]),   .a7(sum30[8]),   .a8(sum30[9]),   .a9(sum30[10]),  .a10(sum30[11]), 
		                .a11(sum30[12]), .a12(sum30[13]), .a13(sum30[14]), .a14(sum30[15]), .a15(sum30[16]), .a16(sum30[17]), .a17(sum30[18]), .a18(sum30[19]), .a19(sum30[20]), .a20(sum30[21]), .a21(sum30[22]),
			        .a22(sum30[23]), .a23(sum30[24]), .a24(sum30[25]), .a25(sum30[26]), .a26(sum30[27]), .a27(sum30[28]), .a28(sum30[29]), .a29(sum30[30]), .a30(sum30[31]), .a31(carry30), 

			        .b0(a[0] & b[31]),   .b1(a[1] & b[31]),   .b2(a[2] & b[31]),   .b3(a[3] & b[31]),   .b4(a[4] & b[31]),   .b5(a[5] & b[31]),   .b6(a[6] & b[31]),   .b7(a[7] & b[31]),
			        .b8(a[8] & b[31]),   .b9(a[9] & b[31]),   .b10(a[10] & b[31]), .b11(a[12] & b[31]), .b12(a[12] & b[31]), .b13(a[13] & b[31]), .b14(a[14] & b[31]), .b15(a[15] & b[31]),
			        .b16(a[16] & b[31]), .b17(a[17] & b[31]), .b18(a[18] & b[31]), .b19(a[19] & b[31]), .b20(a[20] & b[31]), .b21(a[21] & b[31]), .b22(a[22] & b[31]), .b23(a[23] & b[31]),
	                        .b24(a[24] & b[31]), .b25(a[25] & b[31]), .b26(a[26] & b[31]), .b27(a[27] & b[31]), .b28(a[28] & b[31]), .b29(a[29] & b[31]), .b30(a[30] & b[31]), .b31(a[31] & b[31]),	  
	          .cin(1'b0), .cout(carry31));

assign mul[63:1] = {carry31, sum31[31:0], sum30[0], sum29[0], sum28[0], sum27[0], sum26[0], sum25[0], sum24[0], sum23[0], sum22[0], sum21[0], sum20[0], sum19[0], sum18[0], sum17[0], sum16[0], sum15[0], sum14[0], sum13[0], sum12[0], sum11[0], sum10[0], sum9[0], sum8[0], sum7[0], sum6[0], sum5[0], sum4[0], sum3[0], sum2[0], sum1[0]};

endmodule
