module ram (
    input logic clk,
    input logic wr_en,
    input logic [9:0] address,
    input logic [31:0] data_in,
    output logic [31:0] data_out
);

logic [31:0] ram_block [0:1023];

initial begin
    ram_block[0] = 32'b00001_000_0000_0000_0000_00_00111_00000; // R7 mvi
    ram_block[1] = 32'b01110_000_0110_0110_0100_10_00100_10010;
    ram_block[2] = 32'b00000_000_0000_0000_0000_00_01111_00111;
    ram_block[3] = 32'b00001_000_0000_0000_0000_00_10111_00000; // R23 mvi
    ram_block[4] = 32'b11110_110_0110_0110_0110_10_00100_10010;
    ram_block[5] = 32'b00010_000_0000_0000_0000_00_00111_10111; // R7 = R7 + R23
    ram_block[6] = 32'b00011_000_0000_0000_0000_00_10111_00111; // R23 = R23 - R7
    ram_block[7] = 32'b00001_000_0000_0000_0000_00_01000_00000; // R8 mvi
    ram_block[8] = 32'b00000_000_0000_0000_0000_00_11111_11111; // R8 = 1023
    ram_block[9] = 32'b00100_000_0000_0000_0000_00_10010_01000; // ld R18, R8
    ram_block[10] = 32'b00001_000_0000_0000_0000_00_10011_00000; // R19 mvi
    ram_block[11] = 32'b00000_000_0000_0000_0000_00_01101_10110; // 1B6 = 438
    ram_block[12] = 32'b00101_000_0000_0000_0000_00_10010_10011; // st R18, R19
    ram_block[13] = 32'b00000_000_0000_0000_0000_00_00101_10011; // R5 = R19
    ram_block[14] = 32'b00100_000_0000_0000_0000_00_10100_00101; // ld R20, R5
    ram_block[15] = 32'b00110_000_0000_0000_0000_00_10100_00101; // and R20, R5
    ram_block[16] = 32'b00111_000_0000_0000_0000_00_10100_00101; // or R20, R5
    ram_block[17] = 32'b01000_000_0000_0000_0000_00_10100_10010; // xor R20, R18
    ram_block[18] = 32'b01001_000_0000_0000_0000_00_10100_00000; // not R20
    ram_block[1023] = 32'b01110_110_0110_1110_0010_11_00100_10110; // 766E2C96
end

always @(posedge clk) begin
        if(wr_en)
            ram_block[address] <= data_in;
        else
            data_out <= ram_block[address];
end

endmodule
