module multiplexer (
	input logic [31:0] DIN,
	input logic [31:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, R16, R17, R18, R19, R20, R21, R22, R23, R24, R25, R26, R27, R28, R29, R30, R31, G, Sin, Cos,
	input logic R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out, R16out, R17out, R18out, R19out, R20out, R21out, R22out, R23out, R24out, R25out, R26out, R27out, R28out, R29out, R30out, R31out, Gout, DINout, Sinout, Cosout,
	output logic [31:0] BUS
);

logic [35:0] sel;
assign sel [35:0] = {R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out, R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out, R16out, R17out, R18out, R19out, R20out, R21out, R22out, R23out, R24out, R25out, R26out, R27out, R28out, R29out, R30out, R31out, Gout, DINout, Sinout, Cosout};

always @(*) begin
	case (sel) 
		36'b1000_0000_0000_0000_0000_0000_0000_0000_0000: BUS = R0;
		36'b0100_0000_0000_0000_0000_0000_0000_0000_0000: BUS = R1;
		36'b0010_0000_0000_0000_0000_0000_0000_0000_0000: BUS = R2;
		36'b0001_0000_0000_0000_0000_0000_0000_0000_0000: BUS = R3;
		36'b0000_1000_0000_0000_0000_0000_0000_0000_0000: BUS = R4;
		36'b0000_0100_0000_0000_0000_0000_0000_0000_0000: BUS = R5;
		36'b0000_0010_0000_0000_0000_0000_0000_0000_0000: BUS = R6;
		36'b0000_0001_0000_0000_0000_0000_0000_0000_0000: BUS = R7;
		36'b0000_0000_1000_0000_0000_0000_0000_0000_0000: BUS = R8;
		36'b0000_0000_0100_0000_0000_0000_0000_0000_0000: BUS = R9;
		36'b0000_0000_0010_0000_0000_0000_0000_0000_0000: BUS = R10;
		36'b0000_0000_0001_0000_0000_0000_0000_0000_0000: BUS = R11;
		36'b0000_0000_0000_1000_0000_0000_0000_0000_0000: BUS = R12;
		36'b0000_0000_0000_0100_0000_0000_0000_0000_0000: BUS = R13;
		36'b0000_0000_0000_0010_0000_0000_0000_0000_0000: BUS = R14;
		36'b0000_0000_0000_0001_0000_0000_0000_0000_0000: BUS = R15;
		36'b0000_0000_0000_0000_1000_0000_0000_0000_0000: BUS = R16;
		36'b0000_0000_0000_0000_0100_0000_0000_0000_0000: BUS = R17;
		36'b0000_0000_0000_0000_0010_0000_0000_0000_0000: BUS = R18;
		36'b0000_0000_0000_0000_0001_0000_0000_0000_0000: BUS = R19;
		36'b0000_0000_0000_0000_0000_1000_0000_0000_0000: BUS = R20;
		36'b0000_0000_0000_0000_0000_0100_0000_0000_0000: BUS = R21;
		36'b0000_0000_0000_0000_0000_0010_0000_0000_0000: BUS = R22;
		36'b0000_0000_0000_0000_0000_0001_0000_0000_0000: BUS = R23;
		36'b0000_0000_0000_0000_0000_0000_1000_0000_0000: BUS = R24;
		36'b0000_0000_0000_0000_0000_0000_0100_0000_0000: BUS = R25;
		36'b0000_0000_0000_0000_0000_0000_0010_0000_0000: BUS = R26;
		36'b0000_0000_0000_0000_0000_0000_0001_0000_0000: BUS = R27;
		36'b0000_0000_0000_0000_0000_0000_0000_1000_0000: BUS = R28;
		36'b0000_0000_0000_0000_0000_0000_0000_0100_0000: BUS = R29;
		36'b0000_0000_0000_0000_0000_0000_0000_0010_0000: BUS = R30;
		36'b0000_0000_0000_0000_0000_0000_0000_0001_0000: BUS = R31;
		36'b0000_0000_0000_0000_0000_0000_0000_0000_1000: BUS = G;
		36'b0000_0000_0000_0000_0000_0000_0000_0000_0100: BUS = DIN;
		36'b0000_0000_0000_0000_0000_0000_0000_0000_0010: BUS = Sin;
		36'b0000_0000_0000_0000_0000_0000_0000_0000_0001: BUS = Cos;
		default: BUS = 36'b0;
	endcase
end 
endmodule
