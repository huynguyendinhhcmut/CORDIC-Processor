module ram (
    input logic clk,
    input logic wr_en,
    input logic [9:0] address,
    input logic [31:0] data_in,
    output logic [31:0] data_out
);

logic [31:0] ram_block [0:1023];

initial begin
    ram_block[0] = 32'b00001_000_0000_0000_0_00000_00001_00000; // R1 mvi (RX)
    ram_block[1] = 32'b01110_000_0110_0110_0_10010_00100_10010;
    ram_block[2] = 32'b00001_000_0000_0000_0_00000_00010_00000; // R2 mvi
    ram_block[3] = 32'b11110_110_0110_0110_0_11010_00100_10010;
    ram_block[4] = 32'b00010_000_0000_0000_0_00011_00010_00001; // R3 = R1 + R2
    ram_block[5] = 32'b00011_000_0000_0000_0_00100_00011_00010; // R4 = R3 - R2
    ram_block[6] = 32'b00001_000_0000_0000_0_00000_00101_00000; // R5 mvi
    ram_block[7] = 32'b00000_000_0000_0000_0_00000_11111_11111; // R5 = 1023
    ram_block[8] = 32'b00100_000_0000_0000_0_00000_00110_00101; // ld R6, R5
    ram_block[9] = 32'b00001_000_0000_0000_0_00000_00111_00000; // R7 mvi
    ram_block[10] = 32'b00000_000_0000_0000_0_00000_01101_10110; // 1B6 = 438
    ram_block[11] = 32'b00101_000_0000_0000_0_00000_00110_00111; // st R6, R7
    ram_block[12] = 32'b00000_000_0000_0000_0_00000_01000_00111; // R8 = R7
    ram_block[13] = 32'b00100_000_0000_0000_0_00000_01001_01000; // ld R9, R8
    ram_block[14] = 32'b00110_000_0000_0000_0_00000_01001_00101; // and R9, R5
    ram_block[15] = 32'b00111_000_0000_0000_0_00000_01001_00101; // or R9, R5
    ram_block[16] = 32'b01000_000_0000_0000_0_00000_01001_00110; // xor R9, R6
    ram_block[17] = 32'b01001_000_0000_0000_0_00000_01001_00000; // not R9
    ram_block[18] = 32'b00001_000_0000_0000_0_00000_01010_00000; // R10 mvi
    ram_block[19] = 32'b0_10000110_11101100100011100000000; // 246.27734
    ram_block[20] = 32'b00001_000_0000_0000_0_00000_01011_00000; // R11 mvi
    ram_block[21] = 32'b0_10000010_10100110011100011011101; // 13.201383
    ram_block[22] = 32'b10001_000_0000_0000_0_01100_01011_01010; // R12 = R11 + R10
    ram_block[23] = 32'b00001_000_0000_0000_0_00000_01101_00000; // R13 mvi
    ram_block[24] = 32'b0_01111100_11010000101011010010110; // 13 degree
    ram_block[25] = 32'b10100_000_0000_0000_0_00000_01111_01101; // R15 = sin(R13)
    ram_block[26] = 32'b10101_000_0000_0000_0_00000_10000_01101; // R16 = cos(R13)
    ram_block[1023] = 32'b01110_110_0110_1110_0010_11_00100_10110; // 766E2C96
end

always @(posedge clk) begin
        if(wr_en)
            ram_block[address] <= data_in;
        else
            data_out <= ram_block[address];
end

endmodule
