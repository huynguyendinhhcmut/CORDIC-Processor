module multiply32x32 (
	input logic [31:0] a, b,
	output logic [63:0] mul
);

//stage 1
logic [31:0] a1, b1, sum1;
logic cout1;
assign a1[31:0] = {1'b0, (a[31] & b[0]), (a[30] & b[0]), (a[29] & b[0]), (a[28] & b[0]), (a[27] & b[0]), (a[26] & b[0]), (a[25] & b[0]),
					          (a[24] & b[0]), (a[23] & b[0]), (a[22] & b[0]), (a[21] & b[0]), (a[20] & b[0]), (a[19] & b[0]), (a[18] & b[0]), (a[17] & b[0]),
					          (a[16] & b[0]), (a[15] & b[0]), (a[14] & b[0]), (a[13] & b[0]), (a[12] & b[0]), (a[11] & b[0]), (a[10] & b[0]), (a[9] & b[0]),
					          (a[8] & b[0]),  (a[7] & b[0]),  (a[6] & b[0]),  (a[5] & b[0]),  (a[4] & b[0]),  (a[3] & b[0]),  (a[2] & b[0]),  (a[1] & b[0])};
assign b1[31:0] = {(a[31] & b[1]), (a[30] & b[1]), (a[29] & b[1]), (a[28] & b[1]), (a[27] & b[1]), (a[26] & b[1]), (a[25] & b[1]), (a[24] & b[1]), 
						 (a[23] & b[1]), (a[22] & b[1]), (a[21] & b[1]), (a[20] & b[1]), (a[19] & b[1]), (a[18] & b[1]), (a[17] & b[1]), (a[16] & b[1]), 
						 (a[15] & b[1]), (a[14] & b[1]), (a[13] & b[1]), (a[12] & b[1]), (a[11] & b[1]), (a[10] & b[1]), (a[9] & b[1]),  (a[8] & b[1]),  
						 (a[7] & b[1]),  (a[6] & b[1]),  (a[5] & b[1]),  (a[4] & b[1]),  (a[3] & b[1]),  (a[2] & b[1]),  (a[1] & b[1]),  (a[0] & b[1])};
fullAdder32b pa1 (.a(a1), .b(b1), .cin(1'b0), .sum(sum1), .cout(cout1));

//stage2
logic [31:0] a2, b2, sum2;
logic cout2;
assign a2[31:0] = {cout1, sum1[31:1]};
assign b2[31:0] = {(a[31] & b[2]), (a[30] & b[2]), (a[29] & b[2]), (a[28] & b[2]), (a[27] & b[2]), (a[26] & b[2]), (a[25] & b[2]), (a[24] & b[2]), 
						 (a[23] & b[2]), (a[22] & b[2]), (a[21] & b[2]), (a[20] & b[2]), (a[19] & b[2]), (a[18] & b[2]), (a[17] & b[2]), (a[16] & b[2]), 
						 (a[15] & b[2]), (a[14] & b[2]), (a[13] & b[2]), (a[12] & b[2]), (a[11] & b[2]), (a[10] & b[2]), (a[9] & b[2]),  (a[8] & b[2]),  
						 (a[7] & b[2]),  (a[6] & b[2]),  (a[5] & b[2]),  (a[4] & b[2]),  (a[3] & b[2]),  (a[2] & b[2]),  (a[1] & b[2]),  (a[0] & b[2])};
fullAdder32b pa2 (.a(a2), .b(b2), .cin(1'b0), .sum(sum2), .cout(cout2));

//stage3
logic [31:0] a3, b3, sum3;
logic cout3;
assign a3[31:0] = {cout2, sum2[31:1]};
assign b3[31:0] = {(a[31] & b[3]), (a[30] & b[3]), (a[29] & b[3]), (a[28] & b[3]), (a[27] & b[3]), (a[26] & b[3]), (a[25] & b[3]), (a[24] & b[3]), 
						 (a[23] & b[3]), (a[22] & b[3]), (a[21] & b[3]), (a[20] & b[3]), (a[19] & b[3]), (a[18] & b[3]), (a[17] & b[3]), (a[16] & b[3]), 
						 (a[15] & b[3]), (a[14] & b[3]), (a[13] & b[3]), (a[12] & b[3]), (a[11] & b[3]), (a[10] & b[3]), (a[9] & b[3]),  (a[8] & b[3]),  
						 (a[7] & b[3]),  (a[6] & b[3]),  (a[5] & b[3]),  (a[4] & b[3]),  (a[3] & b[3]),  (a[2] & b[3]),  (a[1] & b[3]),  (a[0] & b[3])};
fullAdder32b pa3 (.a(a3), .b(b3), .cin(1'b0), .sum(sum3), .cout(cout3));

//stage4
logic [31:0] a4, b4, sum4;
logic cout4;
assign a4[31:0] = {cout3, sum3[31:1]};
assign b4[31:0] = {(a[31] & b[4]), (a[30] & b[4]), (a[29] & b[4]), (a[28] & b[4]), (a[27] & b[4]), (a[26] & b[4]), (a[25] & b[4]), (a[24] & b[4]), 
						 (a[23] & b[4]), (a[22] & b[4]), (a[21] & b[4]), (a[20] & b[4]), (a[19] & b[4]), (a[18] & b[4]), (a[17] & b[4]), (a[16] & b[4]), 
						 (a[15] & b[4]), (a[14] & b[4]), (a[13] & b[4]), (a[12] & b[4]), (a[11] & b[4]), (a[10] & b[4]), (a[9] & b[4]),  (a[8] & b[4]),  
						 (a[7] & b[4]),  (a[6] & b[4]),  (a[5] & b[4]),  (a[4] & b[4]),  (a[3] & b[4]),  (a[2] & b[4]),  (a[1] & b[4]),  (a[0] & b[4])};
fullAdder32b pa4 (.a(a4), .b(b4), .cin(1'b0), .sum(sum4), .cout(cout4));

//stage5
logic [31:0] a5, b5, sum5;
logic cout5;
assign a5[31:0] = {cout4, sum4[31:1]};
assign b5[31:0] = {(a[31] & b[5]), (a[30] & b[5]), (a[29] & b[5]), (a[28] & b[5]), (a[27] & b[5]), (a[26] & b[5]), (a[25] & b[5]), (a[24] & b[5]), 
						 (a[23] & b[5]), (a[22] & b[5]), (a[21] & b[5]), (a[20] & b[5]), (a[19] & b[5]), (a[18] & b[5]), (a[17] & b[5]), (a[16] & b[5]), 
						 (a[15] & b[5]), (a[14] & b[5]), (a[13] & b[5]), (a[12] & b[5]), (a[11] & b[5]), (a[10] & b[5]), (a[9] & b[5]),  (a[8] & b[5]),  
						 (a[7] & b[5]),  (a[6] & b[5]),  (a[5] & b[5]),  (a[4] & b[5]),  (a[3] & b[5]),  (a[2] & b[5]),  (a[1] & b[5]),  (a[0] & b[5])};
fullAdder32b pa5 (.a(a5), .b(b5), .cin(1'b0), .sum(sum5), .cout(cout5));

//stage6
logic [31:0] a6, b6, sum6;
logic cout6;
assign a6[31:0] = {cout5, sum5[31:1]};
assign b6[31:0] = {(a[31] & b[6]), (a[30] & b[6]), (a[29] & b[6]), (a[28] & b[6]), (a[27] & b[6]), (a[26] & b[6]), (a[25] & b[6]), (a[24] & b[6]), 
						 (a[23] & b[6]), (a[22] & b[6]), (a[21] & b[6]), (a[20] & b[6]), (a[19] & b[6]), (a[18] & b[6]), (a[17] & b[6]), (a[16] & b[6]), 
						 (a[15] & b[6]), (a[14] & b[6]), (a[13] & b[6]), (a[12] & b[6]), (a[11] & b[6]), (a[10] & b[6]), (a[9] & b[6]),  (a[8] & b[6]),  
						 (a[7] & b[6]),  (a[6] & b[6]),  (a[5] & b[6]),  (a[4] & b[6]),  (a[3] & b[6]),  (a[2] & b[6]),  (a[1] & b[6]),  (a[0] & b[6])};
fullAdder32b pa6 (.a(a6), .b(b6), .cin(1'b0), .sum(sum6), .cout(cout6));

//stage7
logic [31:0] a7, b7, sum7;
logic cout7;
assign a7[31:0] = {cout6, sum6[31:1]};
assign b7[31:0] = {(a[31] & b[7]), (a[30] & b[7]), (a[29] & b[7]), (a[28] & b[7]), (a[27] & b[7]), (a[26] & b[7]), (a[25] & b[7]), (a[24] & b[7]), 
						 (a[23] & b[7]), (a[22] & b[7]), (a[21] & b[7]), (a[20] & b[7]), (a[19] & b[7]), (a[18] & b[7]), (a[17] & b[7]), (a[16] & b[7]), 
						 (a[15] & b[7]), (a[14] & b[7]), (a[13] & b[7]), (a[12] & b[7]), (a[11] & b[7]), (a[10] & b[7]), (a[9] & b[7]),  (a[8] & b[7]),  
						 (a[7] & b[7]),  (a[6] & b[7]),  (a[5] & b[7]),  (a[4] & b[7]),  (a[3] & b[7]),  (a[2] & b[7]),  (a[1] & b[7]),  (a[0] & b[7])};
fullAdder32b pa7 (.a(a7), .b(b7), .cin(1'b0), .sum(sum7), .cout(cout7));

//stage8
logic [31:0] a8, b8, sum8;
logic cout8;
assign a8[31:0] = {cout7, sum7[31:1]};
assign b8[31:0] = {(a[31] & b[8]), (a[30] & b[8]), (a[29] & b[8]), (a[28] & b[8]), (a[27] & b[8]), (a[26] & b[8]), (a[25] & b[8]), (a[24] & b[8]), 
						 (a[23] & b[8]), (a[22] & b[8]), (a[21] & b[8]), (a[20] & b[8]), (a[19] & b[8]), (a[18] & b[8]), (a[17] & b[8]), (a[16] & b[8]), 
						 (a[15] & b[8]), (a[14] & b[8]), (a[13] & b[8]), (a[12] & b[8]), (a[11] & b[8]), (a[10] & b[8]), (a[9] & b[8]),  (a[8] & b[8]),  
						 (a[7] & b[8]),  (a[6] & b[8]),  (a[5] & b[8]),  (a[4] & b[8]),  (a[3] & b[8]),  (a[2] & b[8]),  (a[1] & b[8]),  (a[0] & b[8])};
fullAdder32b pa8 (.a(a8), .b(b8), .cin(1'b0), .sum(sum8), .cout(cout8));

//stage9
logic [31:0] a9, b9, sum9;
logic cout9;
assign a9[31:0] = {cout8, sum8[31:1]};
assign b9[31:0] = {(a[31] & b[9]), (a[30] & b[9]), (a[29] & b[9]), (a[28] & b[9]), (a[27] & b[9]), (a[26] & b[9]), (a[25] & b[9]), (a[24] & b[9]), 
						 (a[23] & b[9]), (a[22] & b[9]), (a[21] & b[9]), (a[20] & b[9]), (a[19] & b[9]), (a[18] & b[9]), (a[17] & b[9]), (a[16] & b[9]), 
						 (a[15] & b[9]), (a[14] & b[9]), (a[13] & b[9]), (a[12] & b[9]), (a[11] & b[9]), (a[10] & b[9]), (a[9] & b[9]),  (a[8] & b[9]),  
						 (a[7] & b[9]),  (a[6] & b[9]),  (a[5] & b[9]),  (a[4] & b[9]),  (a[3] & b[9]),  (a[2] & b[9]),  (a[1] & b[9]),  (a[0] & b[9])};
fullAdder32b pa9 (.a(a9), .b(b9), .cin(1'b0), .sum(sum9), .cout(cout9));

//stage10
logic [31:0] a10, b10, sum10;
logic cout10;
assign a10[31:0] = {cout9, sum9[31:1]};
assign b10[31:0] = {(a[31] & b[10]), (a[30] & b[10]), (a[29] & b[10]), (a[28] & b[10]), (a[27] & b[10]), (a[26] & b[10]), (a[25] & b[10]), (a[24] & b[10]), 
						  (a[23] & b[10]), (a[22] & b[10]), (a[21] & b[10]), (a[20] & b[10]), (a[19] & b[10]), (a[18] & b[10]), (a[17] & b[10]), (a[16] & b[10]), 
						  (a[15] & b[10]), (a[14] & b[10]), (a[13] & b[10]), (a[12] & b[10]), (a[11] & b[10]), (a[10] & b[10]), (a[9] & b[10]),  (a[8] & b[10]),  
						  (a[7] & b[10]),  (a[6] & b[10]),  (a[5] & b[10]),  (a[4] & b[10]),  (a[3] & b[10]),  (a[2] & b[10]),  (a[1] & b[10]),  (a[0] & b[10])};
fullAdder32b pa10 (.a(a10), .b(b10), .cin(1'b0), .sum(sum10), .cout(cout10));

//stage11
logic [31:0] a11, b11, sum11;
logic cout11;
assign a11[31:0] = {cout10, sum10[31:1]};
assign b11[31:0] = {(a[31] & b[11]), (a[30] & b[11]), (a[29] & b[11]), (a[28] & b[11]), (a[27] & b[11]), (a[26] & b[11]), (a[25] & b[11]), (a[24] & b[11]), 
						  (a[23] & b[11]), (a[22] & b[11]), (a[21] & b[11]), (a[20] & b[11]), (a[19] & b[11]), (a[18] & b[11]), (a[17] & b[11]), (a[16] & b[11]), 
						  (a[15] & b[11]), (a[14] & b[11]), (a[13] & b[11]), (a[12] & b[11]), (a[11] & b[11]), (a[10] & b[11]), (a[9] & b[11]),  (a[8] & b[11]),  
						  (a[7] & b[11]),  (a[6] & b[11]),  (a[5] & b[11]),  (a[4] & b[11]),  (a[3] & b[11]),  (a[2] & b[11]),  (a[1] & b[11]),  (a[0] & b[11])};
fullAdder32b pa11 (.a(a11), .b(b11), .cin(1'b0), .sum(sum11), .cout(cout11));

//stage12
logic [31:0] a12, b12, sum12;
logic cout12;
assign a12[31:0] = {cout11, sum11[31:1]};
assign b12[31:0] = {(a[31] & b[12]), (a[30] & b[12]), (a[29] & b[12]), (a[28] & b[12]), (a[27] & b[12]), (a[26] & b[12]), (a[25] & b[12]), (a[24] & b[12]), 
						  (a[23] & b[12]), (a[22] & b[12]), (a[21] & b[12]), (a[20] & b[12]), (a[19] & b[12]), (a[18] & b[12]), (a[17] & b[12]), (a[16] & b[12]), 
						  (a[15] & b[12]), (a[14] & b[12]), (a[13] & b[12]), (a[12] & b[12]), (a[11] & b[12]), (a[10] & b[12]), (a[9] & b[12]),  (a[8] & b[12]),  
						  (a[7] & b[12]),  (a[6] & b[12]),  (a[5] & b[12]),  (a[4] & b[12]),  (a[3] & b[12]),  (a[2] & b[12]),  (a[1] & b[12]),  (a[0] & b[12])};
fullAdder32b pa12 (.a(a12), .b(b12), .cin(1'b0), .sum(sum12), .cout(cout12));

//stage13
logic [31:0] a13, b13, sum13;
logic cout13;
assign a13[31:0] = {cout12, sum12[31:1]};
assign b13[31:0] = {(a[31] & b[13]), (a[30] & b[13]), (a[29] & b[13]), (a[28] & b[13]), (a[27] & b[13]), (a[26] & b[13]), (a[25] & b[13]), (a[24] & b[13]), 
						  (a[23] & b[13]), (a[22] & b[13]), (a[21] & b[13]), (a[20] & b[13]), (a[19] & b[13]), (a[18] & b[13]), (a[17] & b[13]), (a[16] & b[13]), 
						  (a[15] & b[13]), (a[14] & b[13]), (a[13] & b[13]), (a[12] & b[13]), (a[11] & b[13]), (a[10] & b[13]), (a[9] & b[13]),  (a[8] & b[13]),  
						  (a[7] & b[13]),  (a[6] & b[13]),  (a[5] & b[13]),  (a[4] & b[13]),  (a[3] & b[13]),  (a[2] & b[13]),  (a[1] & b[13]),  (a[0] & b[13])};
fullAdder32b pa13 (.a(a13), .b(b13), .cin(1'b0), .sum(sum13), .cout(cout13));

//stage14
logic [31:0] a14, b14, sum14;
logic cout14;
assign a14[31:0] = {cout13, sum13[31:1]};
assign b14[31:0] = {(a[31] & b[14]), (a[30] & b[14]), (a[29] & b[14]), (a[28] & b[14]), (a[27] & b[14]), (a[26] & b[14]), (a[25] & b[14]), (a[24] & b[14]), 
						  (a[23] & b[14]), (a[22] & b[14]), (a[21] & b[14]), (a[20] & b[14]), (a[19] & b[14]), (a[18] & b[14]), (a[17] & b[14]), (a[16] & b[14]), 
						  (a[15] & b[14]), (a[14] & b[14]), (a[13] & b[14]), (a[12] & b[14]), (a[11] & b[14]), (a[10] & b[14]), (a[9] & b[14]),  (a[8] & b[14]),  
						  (a[7] & b[14]),  (a[6] & b[14]),  (a[5] & b[14]),  (a[4] & b[14]),  (a[3] & b[14]),  (a[2] & b[14]),  (a[1] & b[14]),  (a[0] & b[14])};
fullAdder32b pa14 (.a(a14), .b(b14), .cin(1'b0), .sum(sum14), .cout(cout14));

//stage15
logic [31:0] a15, b15, sum15;
logic cout15;
assign a15[31:0] = {cout14, sum14[31:1]};
assign b15[31:0] = {(a[31] & b[15]), (a[30] & b[15]), (a[29] & b[15]), (a[28] & b[15]), (a[27] & b[15]), (a[26] & b[15]), (a[25] & b[15]), (a[24] & b[15]), 
						  (a[23] & b[15]), (a[22] & b[15]), (a[21] & b[15]), (a[20] & b[15]), (a[19] & b[15]), (a[18] & b[15]), (a[17] & b[15]), (a[16] & b[15]), 
						  (a[15] & b[15]), (a[14] & b[15]), (a[13] & b[15]), (a[12] & b[15]), (a[11] & b[15]), (a[10] & b[15]), (a[9] & b[15]),  (a[8] & b[15]),  
						  (a[7] & b[15]),  (a[6] & b[15]),  (a[5] & b[15]),  (a[4] & b[15]),  (a[3] & b[15]),  (a[2] & b[15]),  (a[1] & b[15]),  (a[0] & b[15])};
fullAdder32b pa15 (.a(a15), .b(b15), .cin(1'b0), .sum(sum15), .cout(cout15));

//stage16
logic [31:0] a16, b16, sum16;
logic cout16;
assign a16[31:0] = {cout15, sum15[31:1]};
assign b16[31:0] = {(a[31] & b[16]), (a[30] & b[16]), (a[29] & b[16]), (a[28] & b[16]), (a[27] & b[16]), (a[26] & b[16]), (a[25] & b[16]), (a[24] & b[16]), 
						  (a[23] & b[16]), (a[22] & b[16]), (a[21] & b[16]), (a[20] & b[16]), (a[19] & b[16]), (a[18] & b[16]), (a[17] & b[16]), (a[16] & b[16]), 
						  (a[15] & b[16]), (a[14] & b[16]), (a[13] & b[16]), (a[12] & b[16]), (a[11] & b[16]), (a[10] & b[16]), (a[9] & b[16]),  (a[8] & b[16]),  
						  (a[7] & b[16]),  (a[6] & b[16]),  (a[5] & b[16]),  (a[4] & b[16]),  (a[3] & b[16]),  (a[2] & b[16]),  (a[1] & b[16]),  (a[0] & b[16])};
fullAdder32b pa16 (.a(a16), .b(b16), .cin(1'b0), .sum(sum16), .cout(cout16));

//stage17
logic [31:0] a17, b17, sum17;
logic cout17;
assign a17[31:0] = {cout16, sum16[31:1]};
assign b17[31:0] = {(a[31] & b[17]), (a[30] & b[17]), (a[29] & b[17]), (a[28] & b[17]), (a[27] & b[17]), (a[26] & b[17]), (a[25] & b[17]), (a[24] & b[17]), 
						  (a[23] & b[17]), (a[22] & b[17]), (a[21] & b[17]), (a[20] & b[17]), (a[19] & b[17]), (a[18] & b[17]), (a[17] & b[17]), (a[16] & b[17]), 
						  (a[15] & b[17]), (a[14] & b[17]), (a[13] & b[17]), (a[12] & b[17]), (a[11] & b[17]), (a[10] & b[17]), (a[9] & b[17]),  (a[8] & b[17]),  
						  (a[7] & b[17]),  (a[6] & b[17]),  (a[5] & b[17]),  (a[4] & b[17]),  (a[3] & b[17]),  (a[2] & b[17]),  (a[1] & b[17]),  (a[0] & b[17])};
fullAdder32b pa17 (.a(a17), .b(b17), .cin(1'b0), .sum(sum17), .cout(cout17));

//stage18
logic [31:0] a18, b18, sum18;
logic cout18;
assign a18[31:0] = {cout17, sum17[31:1]};
assign b18[31:0] = {(a[31] & b[18]), (a[30] & b[18]), (a[29] & b[18]), (a[28] & b[18]), (a[27] & b[18]), (a[26] & b[18]), (a[25] & b[18]), (a[24] & b[18]), 
						  (a[23] & b[18]), (a[22] & b[18]), (a[21] & b[18]), (a[20] & b[18]), (a[19] & b[18]), (a[18] & b[18]), (a[17] & b[18]), (a[16] & b[18]), 
						  (a[15] & b[18]), (a[14] & b[18]), (a[13] & b[18]), (a[12] & b[18]), (a[11] & b[18]), (a[10] & b[18]), (a[9] & b[18]),  (a[8] & b[18]),  
						  (a[7] & b[18]),  (a[6] & b[18]),  (a[5] & b[18]),  (a[4] & b[18]),  (a[3] & b[18]),  (a[2] & b[18]),  (a[1] & b[18]),  (a[0] & b[18])};
fullAdder32b pa18 (.a(a18), .b(b18), .cin(1'b0), .sum(sum18), .cout(cout18));

//stage19
logic [31:0] a19, b19, sum19;
logic cout19;
assign a19[31:0] = {cout18, sum18[31:1]};
assign b19[31:0] = {(a[31] & b[19]), (a[30] & b[19]), (a[29] & b[19]), (a[28] & b[19]), (a[27] & b[19]), (a[26] & b[19]), (a[25] & b[19]), (a[24] & b[19]), 
						  (a[23] & b[19]), (a[22] & b[19]), (a[21] & b[19]), (a[20] & b[19]), (a[19] & b[19]), (a[18] & b[19]), (a[17] & b[19]), (a[16] & b[19]), 
						  (a[15] & b[19]), (a[14] & b[19]), (a[13] & b[19]), (a[12] & b[19]), (a[11] & b[19]), (a[10] & b[19]), (a[9] & b[19]),  (a[8] & b[19]),  
						  (a[7] & b[19]),  (a[6] & b[19]),  (a[5] & b[19]),  (a[4] & b[19]),  (a[3] & b[19]),  (a[2] & b[19]),  (a[1] & b[19]),  (a[0] & b[19])};
fullAdder32b pa19 (.a(a19), .b(b19), .cin(1'b0), .sum(sum19), .cout(cout19));


//stage20
logic [31:0] a20, b20, sum20;
logic cout20;
assign a20[31:0] = {cout19, sum19[31:1]};
assign b20[31:0] = {(a[31] & b[20]), (a[30] & b[20]), (a[29] & b[20]), (a[28] & b[20]), (a[27] & b[20]), (a[26] & b[20]), (a[25] & b[20]), (a[24] & b[20]), 
						  (a[23] & b[20]), (a[22] & b[20]), (a[21] & b[20]), (a[20] & b[20]), (a[19] & b[20]), (a[18] & b[20]), (a[17] & b[20]), (a[16] & b[20]), 
						  (a[15] & b[20]), (a[14] & b[20]), (a[13] & b[20]), (a[12] & b[20]), (a[11] & b[20]), (a[10] & b[20]), (a[9] & b[20]),  (a[8] & b[20]),  
						  (a[7] & b[20]),  (a[6] & b[20]),  (a[5] & b[20]),  (a[4] & b[20]),  (a[3] & b[20]),  (a[2] & b[20]),  (a[1] & b[20]),  (a[0] & b[20])};
fullAdder32b pa20 (.a(a20), .b(b20), .cin(1'b0), .sum(sum20), .cout(cout20));

//stage21
logic [31:0] a21, b21, sum21;
logic cout21;
assign a21[31:0] = {cout20, sum20[31:1]};
assign b21[31:0] = {(a[31] & b[21]), (a[30] & b[21]), (a[29] & b[21]), (a[28] & b[21]), (a[27] & b[21]), (a[26] & b[21]), (a[25] & b[21]), (a[24] & b[21]), 
						  (a[23] & b[21]), (a[22] & b[21]), (a[21] & b[21]), (a[20] & b[21]), (a[19] & b[21]), (a[18] & b[21]), (a[17] & b[21]), (a[16] & b[21]), 
						  (a[15] & b[21]), (a[14] & b[21]), (a[13] & b[21]), (a[12] & b[21]), (a[11] & b[21]), (a[10] & b[21]), (a[9] & b[21]),  (a[8] & b[21]),  
						  (a[7] & b[21]),  (a[6] & b[21]),  (a[5] & b[21]),  (a[4] & b[21]),  (a[3] & b[21]),  (a[2] & b[21]),  (a[1] & b[21]),  (a[0] & b[21])};
fullAdder32b pa21 (.a(a21), .b(b21), .cin(1'b0), .sum(sum21), .cout(cout21));

//stage22
logic [31:0] a22, b22, sum22;
logic cout22;
assign a22[31:0] = {cout21, sum21[31:1]};
assign b22[31:0] = {(a[31] & b[22]), (a[30] & b[22]), (a[29] & b[22]), (a[28] & b[22]), (a[27] & b[22]), (a[26] & b[22]), (a[25] & b[22]), (a[24] & b[22]), 
						  (a[23] & b[22]), (a[22] & b[22]), (a[21] & b[22]), (a[20] & b[22]), (a[19] & b[22]), (a[18] & b[22]), (a[17] & b[22]), (a[16] & b[22]), 
						  (a[15] & b[22]), (a[14] & b[22]), (a[13] & b[22]), (a[12] & b[22]), (a[11] & b[22]), (a[10] & b[22]), (a[9] & b[22]),  (a[8] & b[22]),  
						  (a[7] & b[22]),  (a[6] & b[22]),  (a[5] & b[22]),  (a[4] & b[22]),  (a[3] & b[22]),  (a[2] & b[22]),  (a[1] & b[22]),  (a[0] & b[22])};
fullAdder32b pa22 (.a(a22), .b(b22), .cin(1'b0), .sum(sum22), .cout(cout22));

//stage23
logic [31:0] a23, b23, sum23;
logic cout23;
assign a23[31:0] = {cout22, sum22[31:1]};
assign b23[31:0] = {(a[31] & b[23]), (a[30] & b[23]), (a[29] & b[23]), (a[28] & b[23]), (a[27] & b[23]), (a[26] & b[23]), (a[25] & b[23]), (a[24] & b[23]), 
						  (a[23] & b[23]), (a[22] & b[23]), (a[21] & b[23]), (a[20] & b[23]), (a[19] & b[23]), (a[18] & b[23]), (a[17] & b[23]), (a[16] & b[23]), 
						  (a[15] & b[23]), (a[14] & b[23]), (a[13] & b[23]), (a[12] & b[23]), (a[11] & b[23]), (a[10] & b[23]), (a[9] & b[23]),  (a[8] & b[23]),  
						  (a[7] & b[23]),  (a[6] & b[23]),  (a[5] & b[23]),  (a[4] & b[23]),  (a[3] & b[23]),  (a[2] & b[23]),  (a[1] & b[23]),  (a[0] & b[23])};
fullAdder32b pa23 (.a(a23), .b(b23), .cin(1'b0), .sum(sum23), .cout(cout23));

//stage24
logic [31:0] a24, b24, sum24;
logic cout24;
assign a24[31:0] = {cout23, sum23[31:1]};
assign b24[31:0] = {(a[31] & b[24]), (a[30] & b[24]), (a[29] & b[24]), (a[28] & b[24]), (a[27] & b[24]), (a[26] & b[24]), (a[25] & b[24]), (a[24] & b[24]), 
						  (a[23] & b[24]), (a[22] & b[24]), (a[21] & b[24]), (a[20] & b[24]), (a[19] & b[24]), (a[18] & b[24]), (a[17] & b[24]), (a[16] & b[24]), 
						  (a[15] & b[24]), (a[14] & b[24]), (a[13] & b[24]), (a[12] & b[24]), (a[11] & b[24]), (a[10] & b[24]), (a[9] & b[24]),  (a[8] & b[24]),  
						  (a[7] & b[24]),  (a[6] & b[24]),  (a[5] & b[24]),  (a[4] & b[24]),  (a[3] & b[24]),  (a[2] & b[24]),  (a[1] & b[24]),  (a[0] & b[24])};
fullAdder32b pa24 (.a(a24), .b(b24), .cin(1'b0), .sum(sum24), .cout(cout24));

//stage25
logic [31:0] a25, b25, sum25;
logic cout25;
assign a25[31:0] = {cout24, sum24[31:1]};
assign b25[31:0] = {(a[31] & b[25]), (a[30] & b[25]), (a[29] & b[25]), (a[28] & b[25]), (a[27] & b[25]), (a[26] & b[25]), (a[25] & b[25]), (a[24] & b[25]), 
						  (a[23] & b[25]), (a[22] & b[25]), (a[21] & b[25]), (a[20] & b[25]), (a[19] & b[25]), (a[18] & b[25]), (a[17] & b[25]), (a[16] & b[25]), 
						  (a[15] & b[25]), (a[14] & b[25]), (a[13] & b[25]), (a[12] & b[25]), (a[11] & b[25]), (a[10] & b[25]), (a[9] & b[25]),  (a[8] & b[25]),  
						  (a[7] & b[25]),  (a[6] & b[25]),  (a[5] & b[25]),  (a[4] & b[25]),  (a[3] & b[25]),  (a[2] & b[25]),  (a[1] & b[25]),  (a[0] & b[25])};
fullAdder32b pa25 (.a(a25), .b(b25), .cin(1'b0), .sum(sum25), .cout(cout25));

//stage26
logic [31:0] a26, b26, sum26;
logic cout26;
assign a26[31:0] = {cout25, sum25[31:1]};
assign b26[31:0] = {(a[31] & b[26]), (a[30] & b[26]), (a[29] & b[26]), (a[28] & b[26]), (a[27] & b[26]), (a[26] & b[26]), (a[25] & b[26]), (a[24] & b[26]), 
						  (a[23] & b[26]), (a[22] & b[26]), (a[21] & b[26]), (a[20] & b[26]), (a[19] & b[26]), (a[18] & b[26]), (a[17] & b[26]), (a[16] & b[26]), 
						  (a[15] & b[26]), (a[14] & b[26]), (a[13] & b[26]), (a[12] & b[26]), (a[11] & b[26]), (a[10] & b[26]), (a[9] & b[26]),  (a[8] & b[26]),  
						  (a[7] & b[26]),  (a[6] & b[26]),  (a[5] & b[26]),  (a[4] & b[26]),  (a[3] & b[26]),  (a[2] & b[26]),  (a[1] & b[26]),  (a[0] & b[26])};
fullAdder32b pa26 (.a(a26), .b(b26), .cin(1'b0), .sum(sum26), .cout(cout26));

//stage27
logic [31:0] a27, b27, sum27;
logic cout27;
assign a27[31:0] = {cout26, sum26[31:1]};
assign b27[31:0] = {(a[31] & b[27]), (a[30] & b[27]), (a[29] & b[27]), (a[28] & b[27]), (a[27] & b[27]), (a[26] & b[27]), (a[25] & b[27]), (a[24] & b[27]), 
						  (a[23] & b[27]), (a[22] & b[27]), (a[21] & b[27]), (a[20] & b[27]), (a[19] & b[27]), (a[18] & b[27]), (a[17] & b[27]), (a[16] & b[27]), 
						  (a[15] & b[27]), (a[14] & b[27]), (a[13] & b[27]), (a[12] & b[27]), (a[11] & b[27]), (a[10] & b[27]), (a[9] & b[27]),  (a[8] & b[27]),  
						  (a[7] & b[27]),  (a[6] & b[27]),  (a[5] & b[27]),  (a[4] & b[27]),  (a[3] & b[27]),  (a[2] & b[27]),  (a[1] & b[27]),  (a[0] & b[27])};
fullAdder32b pa27 (.a(a27), .b(b27), .cin(1'b0), .sum(sum27), .cout(cout27));

//stage28
logic [31:0] a28, b28, sum28;
logic cout28;
assign a28[31:0] = {cout27, sum27[31:1]};
assign b28[31:0] = {(a[31] & b[28]), (a[30] & b[28]), (a[29] & b[28]), (a[28] & b[28]), (a[27] & b[28]), (a[26] & b[28]), (a[25] & b[28]), (a[24] & b[28]), 
						  (a[23] & b[28]), (a[22] & b[28]), (a[21] & b[28]), (a[20] & b[28]), (a[19] & b[28]), (a[18] & b[28]), (a[17] & b[28]), (a[16] & b[28]), 
						  (a[15] & b[28]), (a[14] & b[28]), (a[13] & b[28]), (a[12] & b[28]), (a[11] & b[28]), (a[10] & b[28]), (a[9] & b[28]),  (a[8] & b[28]),  
						  (a[7] & b[28]),  (a[6] & b[28]),  (a[5] & b[28]),  (a[4] & b[28]),  (a[3] & b[28]),  (a[2] & b[28]),  (a[1] & b[28]),  (a[0] & b[28])};
fullAdder32b pa28 (.a(a28), .b(b28), .cin(1'b0), .sum(sum28), .cout(cout28));

//stage29
logic [31:0] a29, b29, sum29;
logic cout29;
assign a29[31:0] = {cout28, sum28[31:1]};
assign b29[31:0] = {(a[31] & b[29]), (a[30] & b[29]), (a[29] & b[29]), (a[28] & b[29]), (a[27] & b[29]), (a[26] & b[29]), (a[25] & b[29]), (a[24] & b[29]), 
						  (a[23] & b[29]), (a[22] & b[29]), (a[21] & b[29]), (a[20] & b[29]), (a[19] & b[29]), (a[18] & b[29]), (a[17] & b[29]), (a[16] & b[29]), 
						  (a[15] & b[29]), (a[14] & b[29]), (a[13] & b[29]), (a[12] & b[29]), (a[11] & b[29]), (a[10] & b[29]), (a[9] & b[29]),  (a[8] & b[29]),  
						  (a[7] & b[29]),  (a[6] & b[29]),  (a[5] & b[29]),  (a[4] & b[29]),  (a[3] & b[29]),  (a[2] & b[29]),  (a[1] & b[29]),  (a[0] & b[29])};
fullAdder32b pa29 (.a(a29), .b(b29), .cin(1'b0), .sum(sum29), .cout(cout29));

//stage30
logic [31:0] a30, b30, sum30;
logic cout30;
assign a30[31:0] = {cout29, sum29[31:1]};
assign b30[31:0] = {(a[31] & b[30]), (a[30] & b[30]), (a[29] & b[30]), (a[28] & b[30]), (a[27] & b[30]), (a[26] & b[30]), (a[25] & b[30]), (a[24] & b[30]), 
						  (a[23] & b[30]), (a[22] & b[30]), (a[21] & b[30]), (a[20] & b[30]), (a[19] & b[30]), (a[18] & b[30]), (a[17] & b[30]), (a[16] & b[30]), 
						  (a[15] & b[30]), (a[14] & b[30]), (a[13] & b[30]), (a[12] & b[30]), (a[11] & b[30]), (a[10] & b[30]), (a[9] & b[30]),  (a[8] & b[30]),  
						  (a[7] & b[30]),  (a[6] & b[30]),  (a[5] & b[30]),  (a[4] & b[30]),  (a[3] & b[30]),  (a[2] & b[30]),  (a[1] & b[30]),  (a[0] & b[30])};
fullAdder32b pa30 (.a(a30), .b(b30), .cin(1'b0), .sum(sum30), .cout(cout30));

//stage31
logic [31:0] a31, b31, sum31;
logic cout31;
assign a31[31:0] = {cout30, sum30[31:1]};
assign b31[31:0] = {(a[31] & b[31]), (a[30] & b[31]), (a[29] & b[31]), (a[28] & b[31]), (a[27] & b[31]), (a[26] & b[31]), (a[25] & b[31]), (a[24] & b[31]), 
						  (a[23] & b[31]), (a[22] & b[31]), (a[21] & b[31]), (a[20] & b[31]), (a[19] & b[31]), (a[18] & b[31]), (a[17] & b[31]), (a[16] & b[31]), 
						  (a[15] & b[31]), (a[14] & b[31]), (a[13] & b[31]), (a[12] & b[31]), (a[11] & b[31]), (a[10] & b[31]), (a[9] & b[31]),  (a[8] & b[31]),  
						  (a[7] & b[31]),  (a[6] & b[31]),  (a[5] & b[31]),  (a[4] & b[31]),  (a[3] & b[31]),  (a[2] & b[31]),  (a[1] & b[31]),  (a[0] & b[31])};
fullAdder32b pa31 (.a(a31), .b(b31), .cin(1'b0), .sum(sum31), .cout(cout31));

assign mul = {cout31,   sum31[31:0], sum30[0], sum29[0], sum28[0], sum27[0], sum26[0], sum25[0], 
				  sum24[0], sum23[0],    sum22[0], sum21[0], sum20[0], sum19[0], sum18[0], sum17[0], 
				  sum16[0], sum15[0],    sum14[0], sum13[0], sum12[0], sum11[0], sum10[0], sum9[0], 
				  sum8[0],  sum7[0],     sum6[0],  sum5[0],  sum4[0],  sum3[0],  sum2[0],  sum1[0], (a[0] & b[0])};

endmodule
